
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f2",x"c4",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"fc",x"f2",x"c4"),
    14 => (x"48",x"e4",x"f9",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f4",x"eb"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"48",x"12",x"1e",x"72"),
    21 => (x"87",x"c4",x"02",x"11"),
    22 => (x"87",x"f6",x"02",x"88"),
    23 => (x"4f",x"26",x"4a",x"26"),
    24 => (x"73",x"1e",x"72",x"1e"),
    25 => (x"11",x"48",x"12",x"1e"),
    26 => (x"4b",x"87",x"ca",x"02"),
    27 => (x"9b",x"98",x"df",x"c3"),
    28 => (x"f0",x"02",x"88",x"73"),
    29 => (x"26",x"4b",x"26",x"87"),
    30 => (x"1e",x"4f",x"26",x"4a"),
    31 => (x"1e",x"72",x"1e",x"73"),
    32 => (x"ca",x"04",x"8b",x"c1"),
    33 => (x"11",x"48",x"12",x"87"),
    34 => (x"88",x"87",x"c4",x"02"),
    35 => (x"26",x"87",x"f1",x"02"),
    36 => (x"26",x"4b",x"26",x"4a"),
    37 => (x"1e",x"74",x"1e",x"4f"),
    38 => (x"1e",x"72",x"1e",x"73"),
    39 => (x"d0",x"04",x"8b",x"c1"),
    40 => (x"11",x"48",x"12",x"87"),
    41 => (x"4c",x"87",x"ca",x"02"),
    42 => (x"9c",x"98",x"df",x"c3"),
    43 => (x"eb",x"02",x"88",x"74"),
    44 => (x"26",x"4a",x"26",x"87"),
    45 => (x"26",x"4c",x"26",x"4b"),
    46 => (x"48",x"73",x"1e",x"4f"),
    47 => (x"02",x"a9",x"73",x"81"),
    48 => (x"53",x"12",x"87",x"c5"),
    49 => (x"26",x"87",x"f6",x"05"),
    50 => (x"66",x"c4",x"1e",x"4f"),
    51 => (x"12",x"48",x"71",x"4a"),
    52 => (x"87",x"fb",x"05",x"51"),
    53 => (x"73",x"1e",x"4f",x"26"),
    54 => (x"a9",x"73",x"81",x"48"),
    55 => (x"f9",x"53",x"72",x"05"),
    56 => (x"0e",x"4f",x"26",x"87"),
    57 => (x"5d",x"5c",x"5b",x"5e"),
    58 => (x"71",x"86",x"f4",x"0e"),
    59 => (x"48",x"a6",x"c4",x"4d"),
    60 => (x"66",x"dc",x"78",x"c0"),
    61 => (x"48",x"a6",x"c8",x"4b"),
    62 => (x"97",x"15",x"78",x"c0"),
    63 => (x"02",x"6e",x"97",x"7e"),
    64 => (x"13",x"87",x"f0",x"c0"),
    65 => (x"da",x"02",x"9c",x"4c"),
    66 => (x"4a",x"6e",x"97",x"87"),
    67 => (x"aa",x"b7",x"49",x"74"),
    68 => (x"c8",x"87",x"c9",x"05"),
    69 => (x"78",x"c1",x"48",x"a6"),
    70 => (x"87",x"c2",x"4c",x"c0"),
    71 => (x"9c",x"74",x"4c",x"13"),
    72 => (x"c8",x"87",x"e6",x"05"),
    73 => (x"87",x"cb",x"02",x"66"),
    74 => (x"c1",x"48",x"66",x"c4"),
    75 => (x"58",x"a6",x"c8",x"80"),
    76 => (x"c4",x"87",x"ff",x"fe"),
    77 => (x"8e",x"f4",x"48",x"66"),
    78 => (x"4c",x"26",x"4d",x"26"),
    79 => (x"4f",x"26",x"4b",x"26"),
    80 => (x"c1",x"4a",x"71",x"1e"),
    81 => (x"04",x"aa",x"b7",x"c1"),
    82 => (x"c6",x"c1",x"87",x"d9"),
    83 => (x"d2",x"01",x"aa",x"b7"),
    84 => (x"48",x"66",x"c4",x"87"),
    85 => (x"ca",x"05",x"a8",x"d0"),
    86 => (x"c0",x"49",x"72",x"87"),
    87 => (x"48",x"71",x"89",x"f7"),
    88 => (x"c1",x"87",x"ec",x"c0"),
    89 => (x"04",x"aa",x"b7",x"e1"),
    90 => (x"e6",x"c1",x"87",x"d8"),
    91 => (x"d1",x"01",x"aa",x"b7"),
    92 => (x"48",x"66",x"c4",x"87"),
    93 => (x"c9",x"05",x"a8",x"d0"),
    94 => (x"c1",x"49",x"72",x"87"),
    95 => (x"48",x"71",x"89",x"d7"),
    96 => (x"f0",x"c0",x"87",x"cd"),
    97 => (x"aa",x"b7",x"c9",x"8a"),
    98 => (x"ff",x"87",x"c2",x"06"),
    99 => (x"26",x"48",x"72",x"4a"),
   100 => (x"5b",x"5e",x"0e",x"4f"),
   101 => (x"f8",x"0e",x"5d",x"5c"),
   102 => (x"c4",x"7e",x"71",x"86"),
   103 => (x"78",x"c0",x"48",x"a6"),
   104 => (x"a7",x"f9",x"c1",x"4c"),
   105 => (x"49",x"66",x"c4",x"1e"),
   106 => (x"c4",x"87",x"f8",x"fc"),
   107 => (x"6e",x"49",x"70",x"86"),
   108 => (x"97",x"83",x"71",x"4b"),
   109 => (x"ed",x"c0",x"49",x"6b"),
   110 => (x"87",x"c6",x"05",x"a9"),
   111 => (x"c1",x"48",x"a6",x"c4"),
   112 => (x"66",x"d8",x"83",x"78"),
   113 => (x"d8",x"87",x"c5",x"02"),
   114 => (x"0b",x"7b",x"0b",x"66"),
   115 => (x"d3",x"05",x"6b",x"97"),
   116 => (x"02",x"66",x"c4",x"87"),
   117 => (x"4a",x"74",x"87",x"c7"),
   118 => (x"c2",x"8a",x"0a",x"c0"),
   119 => (x"72",x"4a",x"74",x"87"),
   120 => (x"87",x"ef",x"c0",x"48"),
   121 => (x"13",x"1e",x"66",x"dc"),
   122 => (x"87",x"d4",x"fd",x"49"),
   123 => (x"4d",x"70",x"86",x"c4"),
   124 => (x"03",x"ad",x"b7",x"c0"),
   125 => (x"66",x"c4",x"87",x"d4"),
   126 => (x"74",x"87",x"c9",x"02"),
   127 => (x"88",x"08",x"c0",x"48"),
   128 => (x"87",x"c2",x"7e",x"70"),
   129 => (x"48",x"6e",x"7e",x"74"),
   130 => (x"66",x"dc",x"87",x"c9"),
   131 => (x"4c",x"a4",x"75",x"94"),
   132 => (x"f8",x"87",x"ef",x"fe"),
   133 => (x"26",x"4d",x"26",x"8e"),
   134 => (x"26",x"4b",x"26",x"4c"),
   135 => (x"1e",x"00",x"20",x"4f"),
   136 => (x"9a",x"72",x"1e",x"73"),
   137 => (x"87",x"e7",x"c0",x"02"),
   138 => (x"4b",x"c1",x"48",x"c0"),
   139 => (x"d1",x"06",x"a9",x"72"),
   140 => (x"06",x"82",x"72",x"87"),
   141 => (x"83",x"73",x"87",x"c9"),
   142 => (x"f4",x"01",x"a9",x"72"),
   143 => (x"c1",x"87",x"c3",x"87"),
   144 => (x"a9",x"72",x"3a",x"b2"),
   145 => (x"80",x"73",x"89",x"03"),
   146 => (x"2b",x"2a",x"c1",x"07"),
   147 => (x"26",x"87",x"f3",x"05"),
   148 => (x"1e",x"4f",x"26",x"4b"),
   149 => (x"4d",x"c4",x"1e",x"75"),
   150 => (x"04",x"a1",x"b7",x"71"),
   151 => (x"81",x"c1",x"b9",x"ff"),
   152 => (x"72",x"07",x"bd",x"c3"),
   153 => (x"ff",x"04",x"a2",x"b7"),
   154 => (x"c1",x"82",x"c1",x"ba"),
   155 => (x"ee",x"fe",x"07",x"bd"),
   156 => (x"04",x"2d",x"c1",x"87"),
   157 => (x"80",x"c1",x"b8",x"ff"),
   158 => (x"ff",x"04",x"2d",x"07"),
   159 => (x"07",x"81",x"c1",x"b9"),
   160 => (x"4f",x"26",x"4d",x"26"),
   161 => (x"ff",x"48",x"11",x"1e"),
   162 => (x"c4",x"78",x"08",x"d4"),
   163 => (x"88",x"c1",x"48",x"66"),
   164 => (x"70",x"58",x"a6",x"c8"),
   165 => (x"87",x"ed",x"05",x"98"),
   166 => (x"ff",x"1e",x"4f",x"26"),
   167 => (x"ff",x"c3",x"48",x"d4"),
   168 => (x"c4",x"51",x"68",x"78"),
   169 => (x"88",x"c1",x"48",x"66"),
   170 => (x"70",x"58",x"a6",x"c8"),
   171 => (x"87",x"eb",x"05",x"98"),
   172 => (x"73",x"1e",x"4f",x"26"),
   173 => (x"4b",x"d4",x"ff",x"1e"),
   174 => (x"6b",x"7b",x"ff",x"c3"),
   175 => (x"7b",x"ff",x"c3",x"4a"),
   176 => (x"32",x"c8",x"49",x"6b"),
   177 => (x"ff",x"c3",x"b1",x"72"),
   178 => (x"c8",x"4a",x"6b",x"7b"),
   179 => (x"c3",x"b2",x"71",x"31"),
   180 => (x"49",x"6b",x"7b",x"ff"),
   181 => (x"b1",x"72",x"32",x"c8"),
   182 => (x"87",x"c4",x"48",x"71"),
   183 => (x"4c",x"26",x"4d",x"26"),
   184 => (x"4f",x"26",x"4b",x"26"),
   185 => (x"5c",x"5b",x"5e",x"0e"),
   186 => (x"4a",x"71",x"0e",x"5d"),
   187 => (x"72",x"4c",x"d4",x"ff"),
   188 => (x"99",x"ff",x"c3",x"49"),
   189 => (x"f9",x"c3",x"7c",x"71"),
   190 => (x"c8",x"05",x"bf",x"e4"),
   191 => (x"48",x"66",x"d0",x"87"),
   192 => (x"a6",x"d4",x"30",x"c9"),
   193 => (x"49",x"66",x"d0",x"58"),
   194 => (x"ff",x"c3",x"29",x"d8"),
   195 => (x"d0",x"7c",x"71",x"99"),
   196 => (x"29",x"d0",x"49",x"66"),
   197 => (x"71",x"99",x"ff",x"c3"),
   198 => (x"49",x"66",x"d0",x"7c"),
   199 => (x"ff",x"c3",x"29",x"c8"),
   200 => (x"d0",x"7c",x"71",x"99"),
   201 => (x"ff",x"c3",x"49",x"66"),
   202 => (x"72",x"7c",x"71",x"99"),
   203 => (x"c3",x"29",x"d0",x"49"),
   204 => (x"7c",x"71",x"99",x"ff"),
   205 => (x"f0",x"c9",x"4b",x"6c"),
   206 => (x"ff",x"c3",x"4d",x"ff"),
   207 => (x"87",x"d0",x"05",x"ab"),
   208 => (x"6c",x"7c",x"ff",x"c3"),
   209 => (x"02",x"8d",x"c1",x"4b"),
   210 => (x"ff",x"c3",x"87",x"c6"),
   211 => (x"87",x"f0",x"02",x"ab"),
   212 => (x"c7",x"fe",x"48",x"73"),
   213 => (x"49",x"c0",x"1e",x"87"),
   214 => (x"c3",x"48",x"d4",x"ff"),
   215 => (x"81",x"c1",x"78",x"ff"),
   216 => (x"a9",x"b7",x"c8",x"c3"),
   217 => (x"26",x"87",x"f1",x"04"),
   218 => (x"1e",x"73",x"1e",x"4f"),
   219 => (x"f8",x"c4",x"87",x"e7"),
   220 => (x"1e",x"c0",x"4b",x"df"),
   221 => (x"c1",x"f0",x"ff",x"c0"),
   222 => (x"e7",x"fd",x"49",x"f7"),
   223 => (x"c1",x"86",x"c4",x"87"),
   224 => (x"ea",x"c0",x"05",x"a8"),
   225 => (x"48",x"d4",x"ff",x"87"),
   226 => (x"c1",x"78",x"ff",x"c3"),
   227 => (x"c0",x"c0",x"c0",x"c0"),
   228 => (x"e1",x"c0",x"1e",x"c0"),
   229 => (x"49",x"e9",x"c1",x"f0"),
   230 => (x"c4",x"87",x"c9",x"fd"),
   231 => (x"05",x"98",x"70",x"86"),
   232 => (x"d4",x"ff",x"87",x"ca"),
   233 => (x"78",x"ff",x"c3",x"48"),
   234 => (x"87",x"cb",x"48",x"c1"),
   235 => (x"c1",x"87",x"e6",x"fe"),
   236 => (x"fd",x"fe",x"05",x"8b"),
   237 => (x"fc",x"48",x"c0",x"87"),
   238 => (x"73",x"1e",x"87",x"e6"),
   239 => (x"48",x"d4",x"ff",x"1e"),
   240 => (x"d3",x"78",x"ff",x"c3"),
   241 => (x"c0",x"1e",x"c0",x"4b"),
   242 => (x"c1",x"c1",x"f0",x"ff"),
   243 => (x"87",x"d4",x"fc",x"49"),
   244 => (x"98",x"70",x"86",x"c4"),
   245 => (x"ff",x"87",x"ca",x"05"),
   246 => (x"ff",x"c3",x"48",x"d4"),
   247 => (x"cb",x"48",x"c1",x"78"),
   248 => (x"87",x"f1",x"fd",x"87"),
   249 => (x"ff",x"05",x"8b",x"c1"),
   250 => (x"48",x"c0",x"87",x"db"),
   251 => (x"0e",x"87",x"f1",x"fb"),
   252 => (x"0e",x"5c",x"5b",x"5e"),
   253 => (x"fd",x"4c",x"d4",x"ff"),
   254 => (x"ea",x"c6",x"87",x"db"),
   255 => (x"f0",x"e1",x"c0",x"1e"),
   256 => (x"fb",x"49",x"c8",x"c1"),
   257 => (x"86",x"c4",x"87",x"de"),
   258 => (x"c8",x"02",x"a8",x"c1"),
   259 => (x"87",x"ea",x"fe",x"87"),
   260 => (x"e2",x"c1",x"48",x"c0"),
   261 => (x"87",x"da",x"fa",x"87"),
   262 => (x"ff",x"cf",x"49",x"70"),
   263 => (x"ea",x"c6",x"99",x"ff"),
   264 => (x"87",x"c8",x"02",x"a9"),
   265 => (x"c0",x"87",x"d3",x"fe"),
   266 => (x"87",x"cb",x"c1",x"48"),
   267 => (x"c0",x"7c",x"ff",x"c3"),
   268 => (x"f4",x"fc",x"4b",x"f1"),
   269 => (x"02",x"98",x"70",x"87"),
   270 => (x"c0",x"87",x"eb",x"c0"),
   271 => (x"f0",x"ff",x"c0",x"1e"),
   272 => (x"fa",x"49",x"fa",x"c1"),
   273 => (x"86",x"c4",x"87",x"de"),
   274 => (x"d9",x"05",x"98",x"70"),
   275 => (x"7c",x"ff",x"c3",x"87"),
   276 => (x"ff",x"c3",x"49",x"6c"),
   277 => (x"7c",x"7c",x"7c",x"7c"),
   278 => (x"02",x"99",x"c0",x"c1"),
   279 => (x"48",x"c1",x"87",x"c4"),
   280 => (x"48",x"c0",x"87",x"d5"),
   281 => (x"ab",x"c2",x"87",x"d1"),
   282 => (x"c0",x"87",x"c4",x"05"),
   283 => (x"c1",x"87",x"c8",x"48"),
   284 => (x"fd",x"fe",x"05",x"8b"),
   285 => (x"f9",x"48",x"c0",x"87"),
   286 => (x"73",x"1e",x"87",x"e4"),
   287 => (x"e4",x"f9",x"c3",x"1e"),
   288 => (x"c7",x"78",x"c1",x"48"),
   289 => (x"48",x"d0",x"ff",x"4b"),
   290 => (x"c8",x"fb",x"78",x"c2"),
   291 => (x"48",x"d0",x"ff",x"87"),
   292 => (x"1e",x"c0",x"78",x"c3"),
   293 => (x"c1",x"d0",x"e5",x"c0"),
   294 => (x"c7",x"f9",x"49",x"c0"),
   295 => (x"c1",x"86",x"c4",x"87"),
   296 => (x"87",x"c1",x"05",x"a8"),
   297 => (x"05",x"ab",x"c2",x"4b"),
   298 => (x"48",x"c0",x"87",x"c5"),
   299 => (x"c1",x"87",x"f9",x"c0"),
   300 => (x"d0",x"ff",x"05",x"8b"),
   301 => (x"87",x"f7",x"fc",x"87"),
   302 => (x"58",x"e8",x"f9",x"c3"),
   303 => (x"cd",x"05",x"98",x"70"),
   304 => (x"c0",x"1e",x"c1",x"87"),
   305 => (x"d0",x"c1",x"f0",x"ff"),
   306 => (x"87",x"d8",x"f8",x"49"),
   307 => (x"d4",x"ff",x"86",x"c4"),
   308 => (x"78",x"ff",x"c3",x"48"),
   309 => (x"c3",x"87",x"e0",x"c4"),
   310 => (x"ff",x"58",x"ec",x"f9"),
   311 => (x"78",x"c2",x"48",x"d0"),
   312 => (x"c3",x"48",x"d4",x"ff"),
   313 => (x"48",x"c1",x"78",x"ff"),
   314 => (x"0e",x"87",x"f5",x"f7"),
   315 => (x"5d",x"5c",x"5b",x"5e"),
   316 => (x"c3",x"4a",x"71",x"0e"),
   317 => (x"d4",x"ff",x"4d",x"ff"),
   318 => (x"ff",x"7c",x"75",x"4c"),
   319 => (x"c3",x"c4",x"48",x"d0"),
   320 => (x"72",x"7c",x"75",x"78"),
   321 => (x"f0",x"ff",x"c0",x"1e"),
   322 => (x"f7",x"49",x"d8",x"c1"),
   323 => (x"86",x"c4",x"87",x"d6"),
   324 => (x"c5",x"02",x"98",x"70"),
   325 => (x"c0",x"48",x"c0",x"87"),
   326 => (x"7c",x"75",x"87",x"f0"),
   327 => (x"c8",x"7c",x"fe",x"c3"),
   328 => (x"66",x"d4",x"1e",x"c0"),
   329 => (x"87",x"dc",x"f5",x"49"),
   330 => (x"7c",x"75",x"86",x"c4"),
   331 => (x"7c",x"75",x"7c",x"75"),
   332 => (x"4b",x"e0",x"da",x"d8"),
   333 => (x"49",x"6c",x"7c",x"75"),
   334 => (x"87",x"c5",x"05",x"99"),
   335 => (x"f3",x"05",x"8b",x"c1"),
   336 => (x"ff",x"7c",x"75",x"87"),
   337 => (x"78",x"c2",x"48",x"d0"),
   338 => (x"cf",x"f6",x"48",x"c1"),
   339 => (x"d4",x"ff",x"1e",x"87"),
   340 => (x"48",x"d0",x"ff",x"4a"),
   341 => (x"c3",x"78",x"d1",x"c4"),
   342 => (x"89",x"c1",x"7a",x"ff"),
   343 => (x"26",x"87",x"f8",x"05"),
   344 => (x"1e",x"73",x"1e",x"4f"),
   345 => (x"ee",x"c5",x"4b",x"71"),
   346 => (x"ff",x"4a",x"df",x"cd"),
   347 => (x"ff",x"c3",x"48",x"d4"),
   348 => (x"c3",x"48",x"68",x"78"),
   349 => (x"c5",x"02",x"a8",x"fe"),
   350 => (x"05",x"8a",x"c1",x"87"),
   351 => (x"9a",x"72",x"87",x"ed"),
   352 => (x"c0",x"87",x"c5",x"05"),
   353 => (x"87",x"ea",x"c0",x"48"),
   354 => (x"cc",x"02",x"9b",x"73"),
   355 => (x"1e",x"66",x"c8",x"87"),
   356 => (x"c5",x"f4",x"49",x"73"),
   357 => (x"c6",x"86",x"c4",x"87"),
   358 => (x"49",x"66",x"c8",x"87"),
   359 => (x"ff",x"87",x"ee",x"fe"),
   360 => (x"ff",x"c3",x"48",x"d4"),
   361 => (x"9b",x"73",x"78",x"78"),
   362 => (x"ff",x"87",x"c5",x"05"),
   363 => (x"78",x"d0",x"48",x"d0"),
   364 => (x"eb",x"f4",x"48",x"c1"),
   365 => (x"1e",x"73",x"1e",x"87"),
   366 => (x"4b",x"c0",x"4a",x"71"),
   367 => (x"c3",x"48",x"d4",x"ff"),
   368 => (x"d0",x"ff",x"78",x"ff"),
   369 => (x"78",x"c3",x"c4",x"48"),
   370 => (x"c3",x"48",x"d4",x"ff"),
   371 => (x"1e",x"72",x"78",x"ff"),
   372 => (x"c1",x"f0",x"ff",x"c0"),
   373 => (x"cb",x"f4",x"49",x"d1"),
   374 => (x"70",x"86",x"c4",x"87"),
   375 => (x"87",x"cd",x"05",x"98"),
   376 => (x"cc",x"1e",x"c0",x"c8"),
   377 => (x"f8",x"fd",x"49",x"66"),
   378 => (x"70",x"86",x"c4",x"87"),
   379 => (x"48",x"d0",x"ff",x"4b"),
   380 => (x"48",x"73",x"78",x"c2"),
   381 => (x"0e",x"87",x"e9",x"f3"),
   382 => (x"5d",x"5c",x"5b",x"5e"),
   383 => (x"c0",x"1e",x"c0",x"0e"),
   384 => (x"c9",x"c1",x"f0",x"ff"),
   385 => (x"87",x"dc",x"f3",x"49"),
   386 => (x"f9",x"c3",x"1e",x"d2"),
   387 => (x"d0",x"fd",x"49",x"ec"),
   388 => (x"c0",x"86",x"c8",x"87"),
   389 => (x"d2",x"84",x"c1",x"4c"),
   390 => (x"f8",x"04",x"ac",x"b7"),
   391 => (x"ec",x"f9",x"c3",x"87"),
   392 => (x"c3",x"49",x"bf",x"97"),
   393 => (x"c0",x"c1",x"99",x"c0"),
   394 => (x"e7",x"c0",x"05",x"a9"),
   395 => (x"f3",x"f9",x"c3",x"87"),
   396 => (x"d0",x"49",x"bf",x"97"),
   397 => (x"f4",x"f9",x"c3",x"31"),
   398 => (x"c8",x"4a",x"bf",x"97"),
   399 => (x"c3",x"b1",x"72",x"32"),
   400 => (x"bf",x"97",x"f5",x"f9"),
   401 => (x"4c",x"71",x"b1",x"4a"),
   402 => (x"ff",x"ff",x"ff",x"cf"),
   403 => (x"ca",x"84",x"c1",x"9c"),
   404 => (x"87",x"e7",x"c1",x"34"),
   405 => (x"97",x"f5",x"f9",x"c3"),
   406 => (x"31",x"c1",x"49",x"bf"),
   407 => (x"f9",x"c3",x"99",x"c6"),
   408 => (x"4a",x"bf",x"97",x"f6"),
   409 => (x"72",x"2a",x"b7",x"c7"),
   410 => (x"f1",x"f9",x"c3",x"b1"),
   411 => (x"4d",x"4a",x"bf",x"97"),
   412 => (x"f9",x"c3",x"9d",x"cf"),
   413 => (x"4a",x"bf",x"97",x"f2"),
   414 => (x"32",x"ca",x"9a",x"c3"),
   415 => (x"97",x"f3",x"f9",x"c3"),
   416 => (x"33",x"c2",x"4b",x"bf"),
   417 => (x"f9",x"c3",x"b2",x"73"),
   418 => (x"4b",x"bf",x"97",x"f4"),
   419 => (x"c6",x"9b",x"c0",x"c3"),
   420 => (x"b2",x"73",x"2b",x"b7"),
   421 => (x"48",x"c1",x"81",x"c2"),
   422 => (x"49",x"70",x"30",x"71"),
   423 => (x"30",x"75",x"48",x"c1"),
   424 => (x"4c",x"72",x"4d",x"70"),
   425 => (x"94",x"71",x"84",x"c1"),
   426 => (x"ad",x"b7",x"c0",x"c8"),
   427 => (x"c1",x"87",x"cc",x"06"),
   428 => (x"c8",x"2d",x"b7",x"34"),
   429 => (x"01",x"ad",x"b7",x"c0"),
   430 => (x"74",x"87",x"f4",x"ff"),
   431 => (x"87",x"dc",x"f0",x"48"),
   432 => (x"5c",x"5b",x"5e",x"0e"),
   433 => (x"86",x"f8",x"0e",x"5d"),
   434 => (x"48",x"d2",x"c2",x"c4"),
   435 => (x"fa",x"c3",x"78",x"c0"),
   436 => (x"49",x"c0",x"1e",x"ca"),
   437 => (x"c4",x"87",x"de",x"fb"),
   438 => (x"05",x"98",x"70",x"86"),
   439 => (x"48",x"c0",x"87",x"c5"),
   440 => (x"c0",x"87",x"ce",x"c9"),
   441 => (x"c0",x"7e",x"c1",x"4d"),
   442 => (x"49",x"bf",x"f9",x"fe"),
   443 => (x"4a",x"c0",x"fb",x"c3"),
   444 => (x"e6",x"4b",x"c8",x"71"),
   445 => (x"98",x"70",x"87",x"c5"),
   446 => (x"c0",x"87",x"c2",x"05"),
   447 => (x"f5",x"fe",x"c0",x"7e"),
   448 => (x"fb",x"c3",x"49",x"bf"),
   449 => (x"c8",x"71",x"4a",x"dc"),
   450 => (x"87",x"ef",x"e5",x"4b"),
   451 => (x"c2",x"05",x"98",x"70"),
   452 => (x"6e",x"7e",x"c0",x"87"),
   453 => (x"87",x"fd",x"c0",x"02"),
   454 => (x"bf",x"d0",x"c1",x"c4"),
   455 => (x"c8",x"c2",x"c4",x"4d"),
   456 => (x"48",x"7e",x"bf",x"9f"),
   457 => (x"a8",x"ea",x"d6",x"c5"),
   458 => (x"c4",x"87",x"c7",x"05"),
   459 => (x"4d",x"bf",x"d0",x"c1"),
   460 => (x"48",x"6e",x"87",x"ce"),
   461 => (x"a8",x"d5",x"e9",x"ca"),
   462 => (x"c0",x"87",x"c5",x"02"),
   463 => (x"87",x"f1",x"c7",x"48"),
   464 => (x"1e",x"ca",x"fa",x"c3"),
   465 => (x"ec",x"f9",x"49",x"75"),
   466 => (x"70",x"86",x"c4",x"87"),
   467 => (x"87",x"c5",x"05",x"98"),
   468 => (x"dc",x"c7",x"48",x"c0"),
   469 => (x"f5",x"fe",x"c0",x"87"),
   470 => (x"fb",x"c3",x"49",x"bf"),
   471 => (x"c8",x"71",x"4a",x"dc"),
   472 => (x"87",x"d7",x"e4",x"4b"),
   473 => (x"c8",x"05",x"98",x"70"),
   474 => (x"d2",x"c2",x"c4",x"87"),
   475 => (x"da",x"78",x"c1",x"48"),
   476 => (x"f9",x"fe",x"c0",x"87"),
   477 => (x"fb",x"c3",x"49",x"bf"),
   478 => (x"c8",x"71",x"4a",x"c0"),
   479 => (x"87",x"fb",x"e3",x"4b"),
   480 => (x"c0",x"02",x"98",x"70"),
   481 => (x"48",x"c0",x"87",x"c5"),
   482 => (x"c4",x"87",x"e6",x"c6"),
   483 => (x"bf",x"97",x"c8",x"c2"),
   484 => (x"a9",x"d5",x"c1",x"49"),
   485 => (x"87",x"cd",x"c0",x"05"),
   486 => (x"97",x"c9",x"c2",x"c4"),
   487 => (x"ea",x"c2",x"49",x"bf"),
   488 => (x"c5",x"c0",x"02",x"a9"),
   489 => (x"c6",x"48",x"c0",x"87"),
   490 => (x"fa",x"c3",x"87",x"c7"),
   491 => (x"7e",x"bf",x"97",x"ca"),
   492 => (x"a8",x"e9",x"c3",x"48"),
   493 => (x"87",x"ce",x"c0",x"02"),
   494 => (x"eb",x"c3",x"48",x"6e"),
   495 => (x"c5",x"c0",x"02",x"a8"),
   496 => (x"c5",x"48",x"c0",x"87"),
   497 => (x"fa",x"c3",x"87",x"eb"),
   498 => (x"49",x"bf",x"97",x"d5"),
   499 => (x"cc",x"c0",x"05",x"99"),
   500 => (x"d6",x"fa",x"c3",x"87"),
   501 => (x"c2",x"49",x"bf",x"97"),
   502 => (x"c5",x"c0",x"02",x"a9"),
   503 => (x"c5",x"48",x"c0",x"87"),
   504 => (x"fa",x"c3",x"87",x"cf"),
   505 => (x"48",x"bf",x"97",x"d7"),
   506 => (x"58",x"ce",x"c2",x"c4"),
   507 => (x"c1",x"48",x"4c",x"70"),
   508 => (x"d2",x"c2",x"c4",x"88"),
   509 => (x"d8",x"fa",x"c3",x"58"),
   510 => (x"75",x"49",x"bf",x"97"),
   511 => (x"d9",x"fa",x"c3",x"81"),
   512 => (x"c8",x"4a",x"bf",x"97"),
   513 => (x"7e",x"a1",x"72",x"32"),
   514 => (x"48",x"df",x"c6",x"c4"),
   515 => (x"fa",x"c3",x"78",x"6e"),
   516 => (x"48",x"bf",x"97",x"da"),
   517 => (x"c4",x"58",x"a6",x"c8"),
   518 => (x"02",x"bf",x"d2",x"c2"),
   519 => (x"c0",x"87",x"d4",x"c2"),
   520 => (x"49",x"bf",x"f5",x"fe"),
   521 => (x"4a",x"dc",x"fb",x"c3"),
   522 => (x"e1",x"4b",x"c8",x"71"),
   523 => (x"98",x"70",x"87",x"cd"),
   524 => (x"87",x"c5",x"c0",x"02"),
   525 => (x"f8",x"c3",x"48",x"c0"),
   526 => (x"ca",x"c2",x"c4",x"87"),
   527 => (x"c6",x"c4",x"4c",x"bf"),
   528 => (x"fa",x"c3",x"5c",x"f3"),
   529 => (x"49",x"bf",x"97",x"ef"),
   530 => (x"fa",x"c3",x"31",x"c8"),
   531 => (x"4a",x"bf",x"97",x"ee"),
   532 => (x"fa",x"c3",x"49",x"a1"),
   533 => (x"4a",x"bf",x"97",x"f0"),
   534 => (x"a1",x"72",x"32",x"d0"),
   535 => (x"f1",x"fa",x"c3",x"49"),
   536 => (x"d8",x"4a",x"bf",x"97"),
   537 => (x"49",x"a1",x"72",x"32"),
   538 => (x"c4",x"91",x"66",x"c4"),
   539 => (x"81",x"bf",x"df",x"c6"),
   540 => (x"59",x"e7",x"c6",x"c4"),
   541 => (x"97",x"f7",x"fa",x"c3"),
   542 => (x"32",x"c8",x"4a",x"bf"),
   543 => (x"97",x"f6",x"fa",x"c3"),
   544 => (x"4a",x"a2",x"4b",x"bf"),
   545 => (x"97",x"f8",x"fa",x"c3"),
   546 => (x"33",x"d0",x"4b",x"bf"),
   547 => (x"c3",x"4a",x"a2",x"73"),
   548 => (x"bf",x"97",x"f9",x"fa"),
   549 => (x"d8",x"9b",x"cf",x"4b"),
   550 => (x"4a",x"a2",x"73",x"33"),
   551 => (x"5a",x"eb",x"c6",x"c4"),
   552 => (x"bf",x"e7",x"c6",x"c4"),
   553 => (x"74",x"8a",x"c2",x"4a"),
   554 => (x"eb",x"c6",x"c4",x"92"),
   555 => (x"78",x"a1",x"72",x"48"),
   556 => (x"c3",x"87",x"ca",x"c1"),
   557 => (x"bf",x"97",x"dc",x"fa"),
   558 => (x"c3",x"31",x"c8",x"49"),
   559 => (x"bf",x"97",x"db",x"fa"),
   560 => (x"c4",x"49",x"a1",x"4a"),
   561 => (x"c4",x"59",x"da",x"c2"),
   562 => (x"49",x"bf",x"d6",x"c2"),
   563 => (x"ff",x"c7",x"31",x"c5"),
   564 => (x"c4",x"29",x"c9",x"81"),
   565 => (x"c3",x"59",x"f3",x"c6"),
   566 => (x"bf",x"97",x"e1",x"fa"),
   567 => (x"c3",x"32",x"c8",x"4a"),
   568 => (x"bf",x"97",x"e0",x"fa"),
   569 => (x"c4",x"4a",x"a2",x"4b"),
   570 => (x"82",x"6e",x"92",x"66"),
   571 => (x"5a",x"ef",x"c6",x"c4"),
   572 => (x"48",x"e7",x"c6",x"c4"),
   573 => (x"c6",x"c4",x"78",x"c0"),
   574 => (x"a1",x"72",x"48",x"e3"),
   575 => (x"f3",x"c6",x"c4",x"78"),
   576 => (x"e7",x"c6",x"c4",x"48"),
   577 => (x"c6",x"c4",x"78",x"bf"),
   578 => (x"c6",x"c4",x"48",x"f7"),
   579 => (x"c4",x"78",x"bf",x"eb"),
   580 => (x"02",x"bf",x"d2",x"c2"),
   581 => (x"74",x"87",x"c9",x"c0"),
   582 => (x"70",x"30",x"c4",x"48"),
   583 => (x"87",x"c9",x"c0",x"7e"),
   584 => (x"bf",x"ef",x"c6",x"c4"),
   585 => (x"70",x"30",x"c4",x"48"),
   586 => (x"d6",x"c2",x"c4",x"7e"),
   587 => (x"c1",x"78",x"6e",x"48"),
   588 => (x"26",x"8e",x"f8",x"48"),
   589 => (x"26",x"4c",x"26",x"4d"),
   590 => (x"0e",x"4f",x"26",x"4b"),
   591 => (x"5d",x"5c",x"5b",x"5e"),
   592 => (x"c4",x"4a",x"71",x"0e"),
   593 => (x"02",x"bf",x"d2",x"c2"),
   594 => (x"4b",x"72",x"87",x"cb"),
   595 => (x"4c",x"72",x"2b",x"c7"),
   596 => (x"c9",x"9c",x"ff",x"c1"),
   597 => (x"c8",x"4b",x"72",x"87"),
   598 => (x"c3",x"4c",x"72",x"2b"),
   599 => (x"c6",x"c4",x"9c",x"ff"),
   600 => (x"c0",x"83",x"bf",x"df"),
   601 => (x"ab",x"bf",x"f1",x"fe"),
   602 => (x"c0",x"87",x"d9",x"02"),
   603 => (x"c3",x"5b",x"f5",x"fe"),
   604 => (x"73",x"1e",x"ca",x"fa"),
   605 => (x"87",x"fd",x"f0",x"49"),
   606 => (x"98",x"70",x"86",x"c4"),
   607 => (x"c0",x"87",x"c5",x"05"),
   608 => (x"87",x"e6",x"c0",x"48"),
   609 => (x"bf",x"d2",x"c2",x"c4"),
   610 => (x"74",x"87",x"d2",x"02"),
   611 => (x"c3",x"91",x"c4",x"49"),
   612 => (x"69",x"81",x"ca",x"fa"),
   613 => (x"ff",x"ff",x"cf",x"4d"),
   614 => (x"cb",x"9d",x"ff",x"ff"),
   615 => (x"c2",x"49",x"74",x"87"),
   616 => (x"ca",x"fa",x"c3",x"91"),
   617 => (x"4d",x"69",x"9f",x"81"),
   618 => (x"c6",x"fe",x"48",x"75"),
   619 => (x"5b",x"5e",x"0e",x"87"),
   620 => (x"1e",x"0e",x"5d",x"5c"),
   621 => (x"1e",x"c0",x"4d",x"71"),
   622 => (x"dc",x"d0",x"49",x"c1"),
   623 => (x"70",x"86",x"c4",x"87"),
   624 => (x"c1",x"02",x"9c",x"4c"),
   625 => (x"c2",x"c4",x"87",x"c2"),
   626 => (x"49",x"75",x"4a",x"da"),
   627 => (x"87",x"d0",x"da",x"ff"),
   628 => (x"c0",x"02",x"98",x"70"),
   629 => (x"4a",x"74",x"87",x"f2"),
   630 => (x"4b",x"cb",x"49",x"75"),
   631 => (x"87",x"f5",x"da",x"ff"),
   632 => (x"c0",x"02",x"98",x"70"),
   633 => (x"1e",x"c0",x"87",x"e2"),
   634 => (x"c7",x"02",x"9c",x"74"),
   635 => (x"48",x"a6",x"c4",x"87"),
   636 => (x"87",x"c5",x"78",x"c0"),
   637 => (x"c1",x"48",x"a6",x"c4"),
   638 => (x"49",x"66",x"c4",x"78"),
   639 => (x"c4",x"87",x"da",x"cf"),
   640 => (x"9c",x"4c",x"70",x"86"),
   641 => (x"87",x"fe",x"fe",x"05"),
   642 => (x"fc",x"26",x"48",x"74"),
   643 => (x"5e",x"0e",x"87",x"e5"),
   644 => (x"0e",x"5d",x"5c",x"5b"),
   645 => (x"9b",x"4b",x"71",x"1e"),
   646 => (x"c0",x"87",x"c5",x"05"),
   647 => (x"87",x"e5",x"c1",x"48"),
   648 => (x"c0",x"4d",x"a3",x"c8"),
   649 => (x"02",x"66",x"d4",x"7d"),
   650 => (x"66",x"d4",x"87",x"c7"),
   651 => (x"c5",x"05",x"bf",x"97"),
   652 => (x"c1",x"48",x"c0",x"87"),
   653 => (x"66",x"d4",x"87",x"cf"),
   654 => (x"87",x"f1",x"fd",x"49"),
   655 => (x"02",x"9c",x"4c",x"70"),
   656 => (x"dc",x"87",x"c0",x"c1"),
   657 => (x"7d",x"69",x"49",x"a4"),
   658 => (x"c4",x"49",x"a4",x"da"),
   659 => (x"69",x"9f",x"4a",x"a3"),
   660 => (x"d2",x"c2",x"c4",x"7a"),
   661 => (x"87",x"d2",x"02",x"bf"),
   662 => (x"9f",x"49",x"a4",x"d4"),
   663 => (x"ff",x"c0",x"49",x"69"),
   664 => (x"48",x"71",x"99",x"ff"),
   665 => (x"7e",x"70",x"30",x"d0"),
   666 => (x"7e",x"c0",x"87",x"c2"),
   667 => (x"6a",x"48",x"49",x"6e"),
   668 => (x"c0",x"7a",x"70",x"80"),
   669 => (x"49",x"a3",x"cc",x"7b"),
   670 => (x"a3",x"d0",x"79",x"6a"),
   671 => (x"74",x"79",x"c0",x"49"),
   672 => (x"c0",x"87",x"c2",x"48"),
   673 => (x"ea",x"fa",x"26",x"48"),
   674 => (x"5b",x"5e",x"0e",x"87"),
   675 => (x"71",x"0e",x"5d",x"5c"),
   676 => (x"f1",x"fe",x"c0",x"4c"),
   677 => (x"74",x"78",x"ff",x"48"),
   678 => (x"ca",x"c1",x"02",x"9c"),
   679 => (x"49",x"a4",x"c8",x"87"),
   680 => (x"c2",x"c1",x"02",x"69"),
   681 => (x"4a",x"66",x"d0",x"87"),
   682 => (x"d4",x"82",x"49",x"6c"),
   683 => (x"66",x"d0",x"5a",x"a6"),
   684 => (x"c2",x"c4",x"b9",x"4d"),
   685 => (x"ff",x"4a",x"bf",x"ce"),
   686 => (x"71",x"99",x"72",x"ba"),
   687 => (x"e4",x"c0",x"02",x"99"),
   688 => (x"4b",x"a4",x"c4",x"87"),
   689 => (x"f2",x"f9",x"49",x"6b"),
   690 => (x"c4",x"7b",x"70",x"87"),
   691 => (x"49",x"bf",x"ca",x"c2"),
   692 => (x"7c",x"71",x"81",x"6c"),
   693 => (x"c2",x"c4",x"b9",x"75"),
   694 => (x"ff",x"4a",x"bf",x"ce"),
   695 => (x"71",x"99",x"72",x"ba"),
   696 => (x"dc",x"ff",x"05",x"99"),
   697 => (x"f9",x"7c",x"75",x"87"),
   698 => (x"73",x"1e",x"87",x"c9"),
   699 => (x"9b",x"4b",x"71",x"1e"),
   700 => (x"c8",x"87",x"c7",x"02"),
   701 => (x"05",x"69",x"49",x"a3"),
   702 => (x"48",x"c0",x"87",x"c5"),
   703 => (x"c4",x"87",x"eb",x"c0"),
   704 => (x"4a",x"bf",x"e3",x"c6"),
   705 => (x"69",x"49",x"a3",x"c4"),
   706 => (x"c4",x"89",x"c2",x"49"),
   707 => (x"91",x"bf",x"ca",x"c2"),
   708 => (x"c4",x"4a",x"a2",x"71"),
   709 => (x"49",x"bf",x"ce",x"c2"),
   710 => (x"a2",x"71",x"99",x"6b"),
   711 => (x"1e",x"66",x"c8",x"4a"),
   712 => (x"d0",x"ea",x"49",x"72"),
   713 => (x"70",x"86",x"c4",x"87"),
   714 => (x"ca",x"f8",x"48",x"49"),
   715 => (x"1e",x"73",x"1e",x"87"),
   716 => (x"02",x"9b",x"4b",x"71"),
   717 => (x"a3",x"c8",x"87",x"c7"),
   718 => (x"c5",x"05",x"69",x"49"),
   719 => (x"c0",x"48",x"c0",x"87"),
   720 => (x"c6",x"c4",x"87",x"eb"),
   721 => (x"c4",x"4a",x"bf",x"e3"),
   722 => (x"49",x"69",x"49",x"a3"),
   723 => (x"c2",x"c4",x"89",x"c2"),
   724 => (x"71",x"91",x"bf",x"ca"),
   725 => (x"c2",x"c4",x"4a",x"a2"),
   726 => (x"6b",x"49",x"bf",x"ce"),
   727 => (x"4a",x"a2",x"71",x"99"),
   728 => (x"72",x"1e",x"66",x"c8"),
   729 => (x"87",x"c3",x"e6",x"49"),
   730 => (x"49",x"70",x"86",x"c4"),
   731 => (x"87",x"c7",x"f7",x"48"),
   732 => (x"5c",x"5b",x"5e",x"0e"),
   733 => (x"71",x"1e",x"0e",x"5d"),
   734 => (x"4c",x"66",x"d4",x"4b"),
   735 => (x"9b",x"73",x"2c",x"c9"),
   736 => (x"87",x"cf",x"c1",x"02"),
   737 => (x"69",x"49",x"a3",x"c8"),
   738 => (x"87",x"c7",x"c1",x"02"),
   739 => (x"d4",x"4d",x"a3",x"d0"),
   740 => (x"c2",x"c4",x"7d",x"66"),
   741 => (x"ff",x"49",x"bf",x"ce"),
   742 => (x"99",x"4a",x"6b",x"b9"),
   743 => (x"03",x"ac",x"71",x"7e"),
   744 => (x"7b",x"c0",x"87",x"cd"),
   745 => (x"4a",x"a3",x"cc",x"7d"),
   746 => (x"6a",x"49",x"a3",x"c4"),
   747 => (x"72",x"87",x"c2",x"79"),
   748 => (x"02",x"9c",x"74",x"8c"),
   749 => (x"1e",x"49",x"87",x"dd"),
   750 => (x"cc",x"fb",x"49",x"73"),
   751 => (x"d4",x"86",x"c4",x"87"),
   752 => (x"ff",x"c7",x"49",x"66"),
   753 => (x"87",x"cb",x"02",x"99"),
   754 => (x"1e",x"ca",x"fa",x"c3"),
   755 => (x"d9",x"fc",x"49",x"73"),
   756 => (x"26",x"86",x"c4",x"87"),
   757 => (x"0e",x"87",x"dc",x"f5"),
   758 => (x"5d",x"5c",x"5b",x"5e"),
   759 => (x"d0",x"86",x"f0",x"0e"),
   760 => (x"e4",x"c0",x"59",x"a6"),
   761 => (x"66",x"cc",x"4b",x"66"),
   762 => (x"48",x"87",x"ca",x"02"),
   763 => (x"7e",x"70",x"80",x"c8"),
   764 => (x"c5",x"05",x"bf",x"6e"),
   765 => (x"c3",x"48",x"c0",x"87"),
   766 => (x"66",x"cc",x"87",x"ec"),
   767 => (x"73",x"84",x"d0",x"4c"),
   768 => (x"48",x"a6",x"c4",x"49"),
   769 => (x"66",x"c4",x"78",x"6c"),
   770 => (x"6e",x"80",x"c4",x"81"),
   771 => (x"66",x"c8",x"78",x"bf"),
   772 => (x"87",x"c6",x"06",x"a9"),
   773 => (x"89",x"66",x"c4",x"49"),
   774 => (x"b7",x"c0",x"4b",x"71"),
   775 => (x"87",x"c4",x"01",x"ab"),
   776 => (x"87",x"c2",x"c3",x"48"),
   777 => (x"c7",x"48",x"66",x"c4"),
   778 => (x"7e",x"70",x"98",x"ff"),
   779 => (x"c9",x"c1",x"02",x"6e"),
   780 => (x"49",x"c0",x"c8",x"87"),
   781 => (x"4a",x"71",x"89",x"6e"),
   782 => (x"4d",x"ca",x"fa",x"c3"),
   783 => (x"b7",x"73",x"85",x"6e"),
   784 => (x"87",x"c1",x"06",x"aa"),
   785 => (x"48",x"49",x"72",x"4a"),
   786 => (x"70",x"80",x"66",x"c4"),
   787 => (x"49",x"8b",x"72",x"7c"),
   788 => (x"99",x"71",x"8a",x"c1"),
   789 => (x"c0",x"87",x"d9",x"02"),
   790 => (x"15",x"48",x"66",x"e0"),
   791 => (x"66",x"e0",x"c0",x"50"),
   792 => (x"c0",x"80",x"c1",x"48"),
   793 => (x"72",x"58",x"a6",x"e4"),
   794 => (x"71",x"8a",x"c1",x"49"),
   795 => (x"87",x"e7",x"05",x"99"),
   796 => (x"66",x"d0",x"1e",x"c1"),
   797 => (x"87",x"d1",x"f8",x"49"),
   798 => (x"b7",x"c0",x"86",x"c4"),
   799 => (x"e3",x"c1",x"06",x"ab"),
   800 => (x"66",x"e0",x"c0",x"87"),
   801 => (x"b7",x"ff",x"c7",x"4d"),
   802 => (x"e2",x"c0",x"06",x"ab"),
   803 => (x"d0",x"1e",x"75",x"87"),
   804 => (x"d5",x"f9",x"49",x"66"),
   805 => (x"85",x"c0",x"c8",x"87"),
   806 => (x"c0",x"c8",x"48",x"6c"),
   807 => (x"c8",x"7c",x"70",x"80"),
   808 => (x"1e",x"c1",x"8b",x"c0"),
   809 => (x"f7",x"49",x"66",x"d4"),
   810 => (x"86",x"c8",x"87",x"df"),
   811 => (x"c3",x"87",x"ee",x"c0"),
   812 => (x"d0",x"1e",x"ca",x"fa"),
   813 => (x"f1",x"f8",x"49",x"66"),
   814 => (x"c3",x"86",x"c4",x"87"),
   815 => (x"73",x"4a",x"ca",x"fa"),
   816 => (x"80",x"6c",x"48",x"49"),
   817 => (x"49",x"73",x"7c",x"70"),
   818 => (x"99",x"71",x"8b",x"c1"),
   819 => (x"12",x"87",x"ce",x"02"),
   820 => (x"85",x"c1",x"7d",x"97"),
   821 => (x"8b",x"c1",x"49",x"73"),
   822 => (x"f2",x"05",x"99",x"71"),
   823 => (x"ab",x"b7",x"c0",x"87"),
   824 => (x"87",x"e1",x"fe",x"01"),
   825 => (x"8e",x"f0",x"48",x"c1"),
   826 => (x"0e",x"87",x"c8",x"f1"),
   827 => (x"5d",x"5c",x"5b",x"5e"),
   828 => (x"9b",x"4b",x"71",x"0e"),
   829 => (x"c8",x"87",x"c7",x"02"),
   830 => (x"05",x"6d",x"4d",x"a3"),
   831 => (x"48",x"ff",x"87",x"c5"),
   832 => (x"d0",x"87",x"fd",x"c0"),
   833 => (x"49",x"6c",x"4c",x"a3"),
   834 => (x"05",x"99",x"ff",x"c7"),
   835 => (x"02",x"6c",x"87",x"d8"),
   836 => (x"1e",x"c1",x"87",x"c9"),
   837 => (x"f0",x"f5",x"49",x"73"),
   838 => (x"c3",x"86",x"c4",x"87"),
   839 => (x"73",x"1e",x"ca",x"fa"),
   840 => (x"87",x"c6",x"f7",x"49"),
   841 => (x"4a",x"6c",x"86",x"c4"),
   842 => (x"c4",x"04",x"aa",x"6d"),
   843 => (x"cf",x"48",x"ff",x"87"),
   844 => (x"7c",x"a2",x"c1",x"87"),
   845 => (x"ff",x"c7",x"49",x"72"),
   846 => (x"ca",x"fa",x"c3",x"99"),
   847 => (x"48",x"69",x"97",x"81"),
   848 => (x"1e",x"87",x"f0",x"ef"),
   849 => (x"4b",x"71",x"1e",x"73"),
   850 => (x"e4",x"c0",x"02",x"9b"),
   851 => (x"f7",x"c6",x"c4",x"87"),
   852 => (x"c2",x"4a",x"73",x"5b"),
   853 => (x"ca",x"c2",x"c4",x"8a"),
   854 => (x"c4",x"92",x"49",x"bf"),
   855 => (x"48",x"bf",x"e3",x"c6"),
   856 => (x"c6",x"c4",x"80",x"72"),
   857 => (x"48",x"71",x"58",x"fb"),
   858 => (x"c2",x"c4",x"30",x"c4"),
   859 => (x"ed",x"c0",x"58",x"da"),
   860 => (x"f3",x"c6",x"c4",x"87"),
   861 => (x"e7",x"c6",x"c4",x"48"),
   862 => (x"c6",x"c4",x"78",x"bf"),
   863 => (x"c6",x"c4",x"48",x"f7"),
   864 => (x"c4",x"78",x"bf",x"eb"),
   865 => (x"02",x"bf",x"d2",x"c2"),
   866 => (x"c2",x"c4",x"87",x"c9"),
   867 => (x"c4",x"49",x"bf",x"ca"),
   868 => (x"c4",x"87",x"c7",x"31"),
   869 => (x"49",x"bf",x"ef",x"c6"),
   870 => (x"c2",x"c4",x"31",x"c4"),
   871 => (x"d6",x"ee",x"59",x"da"),
   872 => (x"5b",x"5e",x"0e",x"87"),
   873 => (x"4a",x"71",x"0e",x"5c"),
   874 => (x"9a",x"72",x"4b",x"c0"),
   875 => (x"87",x"e1",x"c0",x"02"),
   876 => (x"9f",x"49",x"a2",x"da"),
   877 => (x"c2",x"c4",x"4b",x"69"),
   878 => (x"cf",x"02",x"bf",x"d2"),
   879 => (x"49",x"a2",x"d4",x"87"),
   880 => (x"4c",x"49",x"69",x"9f"),
   881 => (x"9c",x"ff",x"ff",x"c0"),
   882 => (x"87",x"c2",x"34",x"d0"),
   883 => (x"49",x"74",x"4c",x"c0"),
   884 => (x"fd",x"49",x"73",x"b3"),
   885 => (x"dc",x"ed",x"87",x"ed"),
   886 => (x"5b",x"5e",x"0e",x"87"),
   887 => (x"f4",x"0e",x"5d",x"5c"),
   888 => (x"c0",x"4a",x"71",x"86"),
   889 => (x"02",x"9a",x"72",x"7e"),
   890 => (x"fa",x"c3",x"87",x"d8"),
   891 => (x"78",x"c0",x"48",x"c6"),
   892 => (x"48",x"fe",x"f9",x"c3"),
   893 => (x"bf",x"f7",x"c6",x"c4"),
   894 => (x"c2",x"fa",x"c3",x"78"),
   895 => (x"f3",x"c6",x"c4",x"48"),
   896 => (x"c2",x"c4",x"78",x"bf"),
   897 => (x"50",x"c0",x"48",x"e7"),
   898 => (x"bf",x"d6",x"c2",x"c4"),
   899 => (x"c6",x"fa",x"c3",x"49"),
   900 => (x"aa",x"71",x"4a",x"bf"),
   901 => (x"87",x"c0",x"c4",x"03"),
   902 => (x"99",x"cf",x"49",x"72"),
   903 => (x"87",x"e1",x"c0",x"05"),
   904 => (x"1e",x"ca",x"fa",x"c3"),
   905 => (x"bf",x"fe",x"f9",x"c3"),
   906 => (x"fe",x"f9",x"c3",x"49"),
   907 => (x"78",x"a1",x"c1",x"48"),
   908 => (x"c0",x"de",x"ff",x"71"),
   909 => (x"c0",x"86",x"c4",x"87"),
   910 => (x"c3",x"48",x"ed",x"fe"),
   911 => (x"cc",x"78",x"ca",x"fa"),
   912 => (x"ed",x"fe",x"c0",x"87"),
   913 => (x"e0",x"c0",x"48",x"bf"),
   914 => (x"f1",x"fe",x"c0",x"80"),
   915 => (x"c6",x"fa",x"c3",x"58"),
   916 => (x"80",x"c1",x"48",x"bf"),
   917 => (x"58",x"ca",x"fa",x"c3"),
   918 => (x"00",x"0f",x"ad",x"27"),
   919 => (x"bf",x"97",x"bf",x"00"),
   920 => (x"c2",x"02",x"9d",x"4d"),
   921 => (x"e5",x"c3",x"87",x"e2"),
   922 => (x"db",x"c2",x"02",x"ad"),
   923 => (x"ed",x"fe",x"c0",x"87"),
   924 => (x"a3",x"cb",x"4b",x"bf"),
   925 => (x"cf",x"4c",x"11",x"49"),
   926 => (x"d2",x"c1",x"05",x"ac"),
   927 => (x"df",x"49",x"75",x"87"),
   928 => (x"cd",x"89",x"c1",x"99"),
   929 => (x"da",x"c2",x"c4",x"91"),
   930 => (x"4a",x"a3",x"c1",x"81"),
   931 => (x"a3",x"c3",x"51",x"12"),
   932 => (x"c5",x"51",x"12",x"4a"),
   933 => (x"51",x"12",x"4a",x"a3"),
   934 => (x"12",x"4a",x"a3",x"c7"),
   935 => (x"4a",x"a3",x"c9",x"51"),
   936 => (x"a3",x"ce",x"51",x"12"),
   937 => (x"d0",x"51",x"12",x"4a"),
   938 => (x"51",x"12",x"4a",x"a3"),
   939 => (x"12",x"4a",x"a3",x"d2"),
   940 => (x"4a",x"a3",x"d4",x"51"),
   941 => (x"a3",x"d6",x"51",x"12"),
   942 => (x"d8",x"51",x"12",x"4a"),
   943 => (x"51",x"12",x"4a",x"a3"),
   944 => (x"12",x"4a",x"a3",x"dc"),
   945 => (x"4a",x"a3",x"de",x"51"),
   946 => (x"7e",x"c1",x"51",x"12"),
   947 => (x"74",x"87",x"f9",x"c0"),
   948 => (x"05",x"99",x"c8",x"49"),
   949 => (x"74",x"87",x"ea",x"c0"),
   950 => (x"05",x"99",x"d0",x"49"),
   951 => (x"66",x"dc",x"87",x"d0"),
   952 => (x"87",x"ca",x"c0",x"02"),
   953 => (x"66",x"dc",x"49",x"73"),
   954 => (x"02",x"98",x"70",x"0f"),
   955 => (x"05",x"6e",x"87",x"d3"),
   956 => (x"c4",x"87",x"c6",x"c0"),
   957 => (x"c0",x"48",x"da",x"c2"),
   958 => (x"ed",x"fe",x"c0",x"50"),
   959 => (x"e7",x"c2",x"48",x"bf"),
   960 => (x"e7",x"c2",x"c4",x"87"),
   961 => (x"7e",x"50",x"c0",x"48"),
   962 => (x"bf",x"d6",x"c2",x"c4"),
   963 => (x"c6",x"fa",x"c3",x"49"),
   964 => (x"aa",x"71",x"4a",x"bf"),
   965 => (x"87",x"c0",x"fc",x"04"),
   966 => (x"bf",x"f7",x"c6",x"c4"),
   967 => (x"87",x"c8",x"c0",x"05"),
   968 => (x"bf",x"d2",x"c2",x"c4"),
   969 => (x"87",x"fe",x"c1",x"02"),
   970 => (x"48",x"f1",x"fe",x"c0"),
   971 => (x"fa",x"c3",x"78",x"ff"),
   972 => (x"e8",x"49",x"bf",x"c2"),
   973 => (x"49",x"70",x"87",x"c5"),
   974 => (x"59",x"c6",x"fa",x"c3"),
   975 => (x"c3",x"48",x"a6",x"c4"),
   976 => (x"78",x"bf",x"c2",x"fa"),
   977 => (x"bf",x"d2",x"c2",x"c4"),
   978 => (x"87",x"d8",x"c0",x"02"),
   979 => (x"cf",x"49",x"66",x"c4"),
   980 => (x"f8",x"ff",x"ff",x"ff"),
   981 => (x"c0",x"02",x"a9",x"99"),
   982 => (x"4d",x"c0",x"87",x"c5"),
   983 => (x"c1",x"87",x"e1",x"c0"),
   984 => (x"87",x"dc",x"c0",x"4d"),
   985 => (x"cf",x"49",x"66",x"c4"),
   986 => (x"a9",x"99",x"f8",x"ff"),
   987 => (x"87",x"c8",x"c0",x"02"),
   988 => (x"c0",x"48",x"a6",x"c8"),
   989 => (x"87",x"c5",x"c0",x"78"),
   990 => (x"c1",x"48",x"a6",x"c8"),
   991 => (x"4d",x"66",x"c8",x"78"),
   992 => (x"c0",x"05",x"9d",x"75"),
   993 => (x"66",x"c4",x"87",x"e0"),
   994 => (x"c4",x"89",x"c2",x"49"),
   995 => (x"4a",x"bf",x"ca",x"c2"),
   996 => (x"e3",x"c6",x"c4",x"91"),
   997 => (x"f9",x"c3",x"4a",x"bf"),
   998 => (x"a1",x"72",x"48",x"fe"),
   999 => (x"c6",x"fa",x"c3",x"78"),
  1000 => (x"f9",x"78",x"c0",x"48"),
  1001 => (x"48",x"c0",x"87",x"e2"),
  1002 => (x"c6",x"e6",x"8e",x"f4"),
  1003 => (x"00",x"00",x"00",x"87"),
  1004 => (x"ff",x"ff",x"ff",x"00"),
  1005 => (x"00",x"0f",x"bd",x"ff"),
  1006 => (x"00",x"0f",x"c6",x"00"),
  1007 => (x"54",x"41",x"46",x"00"),
  1008 => (x"20",x"20",x"32",x"33"),
  1009 => (x"41",x"46",x"00",x"20"),
  1010 => (x"20",x"36",x"31",x"54"),
  1011 => (x"1e",x"00",x"20",x"20"),
  1012 => (x"c3",x"48",x"d4",x"ff"),
  1013 => (x"48",x"68",x"78",x"ff"),
  1014 => (x"ff",x"1e",x"4f",x"26"),
  1015 => (x"ff",x"c3",x"48",x"d4"),
  1016 => (x"48",x"d0",x"ff",x"78"),
  1017 => (x"ff",x"78",x"e1",x"c8"),
  1018 => (x"78",x"d4",x"48",x"d4"),
  1019 => (x"48",x"fb",x"c6",x"c4"),
  1020 => (x"50",x"bf",x"d4",x"ff"),
  1021 => (x"ff",x"1e",x"4f",x"26"),
  1022 => (x"e0",x"c0",x"48",x"d0"),
  1023 => (x"1e",x"4f",x"26",x"78"),
  1024 => (x"70",x"87",x"cc",x"ff"),
  1025 => (x"c6",x"02",x"99",x"49"),
  1026 => (x"a9",x"fb",x"c0",x"87"),
  1027 => (x"71",x"87",x"f1",x"05"),
  1028 => (x"0e",x"4f",x"26",x"48"),
  1029 => (x"0e",x"5c",x"5b",x"5e"),
  1030 => (x"4c",x"c0",x"4b",x"71"),
  1031 => (x"70",x"87",x"f0",x"fe"),
  1032 => (x"c0",x"02",x"99",x"49"),
  1033 => (x"ec",x"c0",x"87",x"f9"),
  1034 => (x"f2",x"c0",x"02",x"a9"),
  1035 => (x"a9",x"fb",x"c0",x"87"),
  1036 => (x"87",x"eb",x"c0",x"02"),
  1037 => (x"ac",x"b7",x"66",x"cc"),
  1038 => (x"d0",x"87",x"c7",x"03"),
  1039 => (x"87",x"c2",x"02",x"66"),
  1040 => (x"99",x"71",x"53",x"71"),
  1041 => (x"c1",x"87",x"c2",x"02"),
  1042 => (x"87",x"c3",x"fe",x"84"),
  1043 => (x"02",x"99",x"49",x"70"),
  1044 => (x"ec",x"c0",x"87",x"cd"),
  1045 => (x"87",x"c7",x"02",x"a9"),
  1046 => (x"05",x"a9",x"fb",x"c0"),
  1047 => (x"d0",x"87",x"d5",x"ff"),
  1048 => (x"87",x"c3",x"02",x"66"),
  1049 => (x"c0",x"7b",x"97",x"c0"),
  1050 => (x"c4",x"05",x"a9",x"ec"),
  1051 => (x"c5",x"4a",x"74",x"87"),
  1052 => (x"c0",x"4a",x"74",x"87"),
  1053 => (x"48",x"72",x"8a",x"0a"),
  1054 => (x"4d",x"26",x"87",x"c2"),
  1055 => (x"4b",x"26",x"4c",x"26"),
  1056 => (x"fd",x"1e",x"4f",x"26"),
  1057 => (x"49",x"70",x"87",x"c9"),
  1058 => (x"a9",x"b7",x"f0",x"c0"),
  1059 => (x"c0",x"87",x"ca",x"04"),
  1060 => (x"01",x"a9",x"b7",x"f9"),
  1061 => (x"f0",x"c0",x"87",x"c3"),
  1062 => (x"b7",x"c1",x"c1",x"89"),
  1063 => (x"87",x"ca",x"04",x"a9"),
  1064 => (x"a9",x"b7",x"da",x"c1"),
  1065 => (x"c0",x"87",x"c3",x"01"),
  1066 => (x"48",x"71",x"89",x"f7"),
  1067 => (x"5e",x"0e",x"4f",x"26"),
  1068 => (x"71",x"0e",x"5c",x"5b"),
  1069 => (x"4c",x"d4",x"ff",x"4a"),
  1070 => (x"ea",x"c0",x"49",x"72"),
  1071 => (x"9b",x"4b",x"70",x"87"),
  1072 => (x"c1",x"87",x"c2",x"02"),
  1073 => (x"48",x"d0",x"ff",x"8b"),
  1074 => (x"c1",x"78",x"c5",x"c8"),
  1075 => (x"49",x"73",x"7c",x"d5"),
  1076 => (x"f7",x"c3",x"31",x"c6"),
  1077 => (x"4a",x"bf",x"97",x"fc"),
  1078 => (x"70",x"b0",x"71",x"48"),
  1079 => (x"48",x"d0",x"ff",x"7c"),
  1080 => (x"48",x"73",x"78",x"c4"),
  1081 => (x"0e",x"87",x"d5",x"fe"),
  1082 => (x"5d",x"5c",x"5b",x"5e"),
  1083 => (x"71",x"86",x"f8",x"0e"),
  1084 => (x"fb",x"7e",x"c0",x"4c"),
  1085 => (x"4b",x"c0",x"87",x"e4"),
  1086 => (x"97",x"d4",x"c6",x"c1"),
  1087 => (x"a9",x"c0",x"49",x"bf"),
  1088 => (x"fb",x"87",x"cf",x"04"),
  1089 => (x"83",x"c1",x"87",x"f9"),
  1090 => (x"97",x"d4",x"c6",x"c1"),
  1091 => (x"06",x"ab",x"49",x"bf"),
  1092 => (x"c6",x"c1",x"87",x"f1"),
  1093 => (x"02",x"bf",x"97",x"d4"),
  1094 => (x"f2",x"fa",x"87",x"cf"),
  1095 => (x"99",x"49",x"70",x"87"),
  1096 => (x"c0",x"87",x"c6",x"02"),
  1097 => (x"f1",x"05",x"a9",x"ec"),
  1098 => (x"fa",x"4b",x"c0",x"87"),
  1099 => (x"4d",x"70",x"87",x"e1"),
  1100 => (x"c8",x"87",x"dc",x"fa"),
  1101 => (x"d6",x"fa",x"58",x"a6"),
  1102 => (x"c1",x"4a",x"70",x"87"),
  1103 => (x"49",x"a4",x"c8",x"83"),
  1104 => (x"ad",x"49",x"69",x"97"),
  1105 => (x"c0",x"87",x"c7",x"02"),
  1106 => (x"c0",x"05",x"ad",x"ff"),
  1107 => (x"a4",x"c9",x"87",x"e7"),
  1108 => (x"49",x"69",x"97",x"49"),
  1109 => (x"02",x"a9",x"66",x"c4"),
  1110 => (x"c0",x"48",x"87",x"c7"),
  1111 => (x"d4",x"05",x"a8",x"ff"),
  1112 => (x"49",x"a4",x"ca",x"87"),
  1113 => (x"aa",x"49",x"69",x"97"),
  1114 => (x"c0",x"87",x"c6",x"02"),
  1115 => (x"c4",x"05",x"aa",x"ff"),
  1116 => (x"d0",x"7e",x"c1",x"87"),
  1117 => (x"ad",x"ec",x"c0",x"87"),
  1118 => (x"c0",x"87",x"c6",x"02"),
  1119 => (x"c4",x"05",x"ad",x"fb"),
  1120 => (x"c1",x"4b",x"c0",x"87"),
  1121 => (x"fe",x"02",x"6e",x"7e"),
  1122 => (x"e9",x"f9",x"87",x"e1"),
  1123 => (x"f8",x"48",x"73",x"87"),
  1124 => (x"87",x"e6",x"fb",x"8e"),
  1125 => (x"5b",x"5e",x"0e",x"00"),
  1126 => (x"1e",x"0e",x"5d",x"5c"),
  1127 => (x"4c",x"c0",x"4b",x"71"),
  1128 => (x"c0",x"04",x"ab",x"4d"),
  1129 => (x"c3",x"c1",x"87",x"e8"),
  1130 => (x"9d",x"75",x"1e",x"e7"),
  1131 => (x"c0",x"87",x"c4",x"02"),
  1132 => (x"c1",x"87",x"c2",x"4a"),
  1133 => (x"f0",x"49",x"72",x"4a"),
  1134 => (x"86",x"c4",x"87",x"df"),
  1135 => (x"84",x"c1",x"7e",x"70"),
  1136 => (x"87",x"c2",x"05",x"6e"),
  1137 => (x"85",x"c1",x"4c",x"73"),
  1138 => (x"ff",x"06",x"ac",x"73"),
  1139 => (x"48",x"6e",x"87",x"d8"),
  1140 => (x"26",x"4d",x"26",x"26"),
  1141 => (x"26",x"4b",x"26",x"4c"),
  1142 => (x"4a",x"71",x"1e",x"4f"),
  1143 => (x"99",x"ff",x"c3",x"49"),
  1144 => (x"71",x"48",x"d4",x"ff"),
  1145 => (x"c8",x"49",x"72",x"78"),
  1146 => (x"ff",x"c3",x"29",x"b7"),
  1147 => (x"72",x"78",x"71",x"99"),
  1148 => (x"29",x"b7",x"d0",x"49"),
  1149 => (x"71",x"99",x"ff",x"c3"),
  1150 => (x"d8",x"49",x"72",x"78"),
  1151 => (x"ff",x"c3",x"29",x"b7"),
  1152 => (x"26",x"78",x"71",x"99"),
  1153 => (x"5b",x"5e",x"0e",x"4f"),
  1154 => (x"1e",x"0e",x"5d",x"5c"),
  1155 => (x"4b",x"c0",x"4a",x"71"),
  1156 => (x"e3",x"c1",x"49",x"72"),
  1157 => (x"98",x"70",x"87",x"d6"),
  1158 => (x"c1",x"87",x"da",x"05"),
  1159 => (x"c1",x"49",x"74",x"4c"),
  1160 => (x"70",x"87",x"e3",x"e4"),
  1161 => (x"87",x"c2",x"05",x"98"),
  1162 => (x"84",x"c1",x"4b",x"c1"),
  1163 => (x"bf",x"de",x"cb",x"c4"),
  1164 => (x"e8",x"06",x"ac",x"b7"),
  1165 => (x"48",x"d0",x"ff",x"87"),
  1166 => (x"ff",x"78",x"e1",x"c8"),
  1167 => (x"78",x"dd",x"48",x"d4"),
  1168 => (x"c7",x"02",x"9b",x"73"),
  1169 => (x"c6",x"cc",x"c4",x"87"),
  1170 => (x"87",x"c2",x"4d",x"bf"),
  1171 => (x"49",x"75",x"4d",x"c0"),
  1172 => (x"73",x"87",x"c6",x"fe"),
  1173 => (x"87",x"c7",x"02",x"9b"),
  1174 => (x"bf",x"c6",x"cc",x"c4"),
  1175 => (x"c0",x"87",x"c2",x"7e"),
  1176 => (x"fd",x"49",x"6e",x"7e"),
  1177 => (x"49",x"c0",x"87",x"f3"),
  1178 => (x"c0",x"87",x"ee",x"fd"),
  1179 => (x"87",x"e9",x"fd",x"49"),
  1180 => (x"c0",x"48",x"d0",x"ff"),
  1181 => (x"1e",x"c1",x"78",x"e0"),
  1182 => (x"f2",x"c0",x"49",x"dc"),
  1183 => (x"48",x"73",x"87",x"db"),
  1184 => (x"cc",x"fd",x"8e",x"f8"),
  1185 => (x"5b",x"5e",x"0e",x"87"),
  1186 => (x"1e",x"0e",x"5d",x"5c"),
  1187 => (x"de",x"49",x"4c",x"71"),
  1188 => (x"d5",x"c7",x"c4",x"91"),
  1189 => (x"97",x"85",x"71",x"4d"),
  1190 => (x"dd",x"c1",x"02",x"6d"),
  1191 => (x"c0",x"c7",x"c4",x"87"),
  1192 => (x"82",x"74",x"4a",x"bf"),
  1193 => (x"ec",x"fb",x"49",x"72"),
  1194 => (x"6e",x"7e",x"70",x"87"),
  1195 => (x"87",x"f3",x"c0",x"02"),
  1196 => (x"4b",x"c8",x"c7",x"c4"),
  1197 => (x"49",x"cb",x"4a",x"6e"),
  1198 => (x"87",x"fd",x"f7",x"fe"),
  1199 => (x"93",x"cb",x"4b",x"74"),
  1200 => (x"83",x"e4",x"ed",x"c1"),
  1201 => (x"cb",x"c1",x"83",x"c4"),
  1202 => (x"49",x"74",x"7b",x"fe"),
  1203 => (x"87",x"ff",x"c4",x"c1"),
  1204 => (x"c7",x"c4",x"7b",x"75"),
  1205 => (x"49",x"bf",x"97",x"d4"),
  1206 => (x"c8",x"c7",x"c4",x"1e"),
  1207 => (x"d0",x"eb",x"c2",x"49"),
  1208 => (x"74",x"86",x"c4",x"87"),
  1209 => (x"e6",x"c4",x"c1",x"49"),
  1210 => (x"c1",x"49",x"c0",x"87"),
  1211 => (x"c4",x"87",x"c5",x"c6"),
  1212 => (x"c0",x"48",x"fc",x"c6"),
  1213 => (x"dd",x"49",x"c1",x"78"),
  1214 => (x"fb",x"26",x"87",x"d2"),
  1215 => (x"6f",x"4c",x"87",x"d3"),
  1216 => (x"6e",x"69",x"64",x"61"),
  1217 => (x"2e",x"2e",x"2e",x"67"),
  1218 => (x"5b",x"5e",x"0e",x"00"),
  1219 => (x"4b",x"71",x"0e",x"5c"),
  1220 => (x"c0",x"c7",x"c4",x"4a"),
  1221 => (x"49",x"72",x"82",x"bf"),
  1222 => (x"70",x"87",x"fa",x"f9"),
  1223 => (x"c4",x"02",x"9c",x"4c"),
  1224 => (x"fc",x"e9",x"49",x"87"),
  1225 => (x"c0",x"c7",x"c4",x"87"),
  1226 => (x"c1",x"78",x"c0",x"48"),
  1227 => (x"87",x"dc",x"dc",x"49"),
  1228 => (x"0e",x"87",x"e0",x"fa"),
  1229 => (x"5d",x"5c",x"5b",x"5e"),
  1230 => (x"c3",x"86",x"f4",x"0e"),
  1231 => (x"c0",x"4d",x"ca",x"fa"),
  1232 => (x"48",x"a6",x"c4",x"4c"),
  1233 => (x"c7",x"c4",x"78",x"c0"),
  1234 => (x"c0",x"49",x"bf",x"c0"),
  1235 => (x"c1",x"c1",x"06",x"a9"),
  1236 => (x"ca",x"fa",x"c3",x"87"),
  1237 => (x"c0",x"02",x"98",x"48"),
  1238 => (x"c3",x"c1",x"87",x"f8"),
  1239 => (x"66",x"c8",x"1e",x"e7"),
  1240 => (x"c4",x"87",x"c7",x"02"),
  1241 => (x"78",x"c0",x"48",x"a6"),
  1242 => (x"a6",x"c4",x"87",x"c5"),
  1243 => (x"c4",x"78",x"c1",x"48"),
  1244 => (x"e4",x"e9",x"49",x"66"),
  1245 => (x"70",x"86",x"c4",x"87"),
  1246 => (x"c4",x"84",x"c1",x"4d"),
  1247 => (x"80",x"c1",x"48",x"66"),
  1248 => (x"c4",x"58",x"a6",x"c8"),
  1249 => (x"49",x"bf",x"c0",x"c7"),
  1250 => (x"87",x"c6",x"03",x"ac"),
  1251 => (x"ff",x"05",x"9d",x"75"),
  1252 => (x"4c",x"c0",x"87",x"c8"),
  1253 => (x"c3",x"02",x"9d",x"75"),
  1254 => (x"c3",x"c1",x"87",x"e0"),
  1255 => (x"66",x"c8",x"1e",x"e7"),
  1256 => (x"cc",x"87",x"c7",x"02"),
  1257 => (x"78",x"c0",x"48",x"a6"),
  1258 => (x"a6",x"cc",x"87",x"c5"),
  1259 => (x"cc",x"78",x"c1",x"48"),
  1260 => (x"e4",x"e8",x"49",x"66"),
  1261 => (x"70",x"86",x"c4",x"87"),
  1262 => (x"c2",x"02",x"6e",x"7e"),
  1263 => (x"49",x"6e",x"87",x"e9"),
  1264 => (x"69",x"97",x"81",x"cb"),
  1265 => (x"02",x"99",x"d0",x"49"),
  1266 => (x"c1",x"87",x"d6",x"c1"),
  1267 => (x"74",x"4a",x"c9",x"cc"),
  1268 => (x"c1",x"91",x"cb",x"49"),
  1269 => (x"72",x"81",x"e4",x"ed"),
  1270 => (x"c3",x"81",x"c8",x"79"),
  1271 => (x"49",x"74",x"51",x"ff"),
  1272 => (x"c7",x"c4",x"91",x"de"),
  1273 => (x"85",x"71",x"4d",x"d5"),
  1274 => (x"7d",x"97",x"c1",x"c2"),
  1275 => (x"c0",x"49",x"a5",x"c1"),
  1276 => (x"c2",x"c4",x"51",x"e0"),
  1277 => (x"02",x"bf",x"97",x"da"),
  1278 => (x"84",x"c1",x"87",x"d2"),
  1279 => (x"c4",x"4b",x"a5",x"c2"),
  1280 => (x"db",x"4a",x"da",x"c2"),
  1281 => (x"f0",x"f2",x"fe",x"49"),
  1282 => (x"87",x"db",x"c1",x"87"),
  1283 => (x"c0",x"49",x"a5",x"cd"),
  1284 => (x"c2",x"84",x"c1",x"51"),
  1285 => (x"4a",x"6e",x"4b",x"a5"),
  1286 => (x"f2",x"fe",x"49",x"cb"),
  1287 => (x"c6",x"c1",x"87",x"db"),
  1288 => (x"c5",x"ca",x"c1",x"87"),
  1289 => (x"cb",x"49",x"74",x"4a"),
  1290 => (x"e4",x"ed",x"c1",x"91"),
  1291 => (x"c4",x"79",x"72",x"81"),
  1292 => (x"bf",x"97",x"da",x"c2"),
  1293 => (x"74",x"87",x"d8",x"02"),
  1294 => (x"c1",x"91",x"de",x"49"),
  1295 => (x"d5",x"c7",x"c4",x"84"),
  1296 => (x"c4",x"83",x"71",x"4b"),
  1297 => (x"dd",x"4a",x"da",x"c2"),
  1298 => (x"ec",x"f1",x"fe",x"49"),
  1299 => (x"74",x"87",x"d8",x"87"),
  1300 => (x"c4",x"93",x"de",x"4b"),
  1301 => (x"cb",x"83",x"d5",x"c7"),
  1302 => (x"51",x"c0",x"49",x"a3"),
  1303 => (x"6e",x"73",x"84",x"c1"),
  1304 => (x"fe",x"49",x"cb",x"4a"),
  1305 => (x"c4",x"87",x"d2",x"f1"),
  1306 => (x"80",x"c1",x"48",x"66"),
  1307 => (x"c7",x"58",x"a6",x"c8"),
  1308 => (x"c5",x"c0",x"03",x"ac"),
  1309 => (x"fc",x"05",x"6e",x"87"),
  1310 => (x"48",x"74",x"87",x"e0"),
  1311 => (x"d0",x"f5",x"8e",x"f4"),
  1312 => (x"1e",x"73",x"1e",x"87"),
  1313 => (x"cb",x"49",x"4b",x"71"),
  1314 => (x"e4",x"ed",x"c1",x"91"),
  1315 => (x"4a",x"a1",x"c8",x"81"),
  1316 => (x"48",x"fc",x"f7",x"c3"),
  1317 => (x"a1",x"c9",x"50",x"12"),
  1318 => (x"d4",x"c6",x"c1",x"4a"),
  1319 => (x"ca",x"50",x"12",x"48"),
  1320 => (x"d4",x"c7",x"c4",x"81"),
  1321 => (x"c4",x"50",x"11",x"48"),
  1322 => (x"bf",x"97",x"d4",x"c7"),
  1323 => (x"49",x"c0",x"1e",x"49"),
  1324 => (x"87",x"fd",x"e3",x"c2"),
  1325 => (x"48",x"fc",x"c6",x"c4"),
  1326 => (x"49",x"c1",x"78",x"de"),
  1327 => (x"26",x"87",x"cd",x"d6"),
  1328 => (x"1e",x"87",x"d2",x"f4"),
  1329 => (x"cb",x"49",x"4a",x"71"),
  1330 => (x"e4",x"ed",x"c1",x"91"),
  1331 => (x"11",x"81",x"c8",x"81"),
  1332 => (x"c0",x"c7",x"c4",x"48"),
  1333 => (x"c0",x"c7",x"c4",x"58"),
  1334 => (x"c1",x"78",x"c0",x"48"),
  1335 => (x"87",x"ec",x"d5",x"49"),
  1336 => (x"c0",x"1e",x"4f",x"26"),
  1337 => (x"cb",x"fe",x"c0",x"49"),
  1338 => (x"1e",x"4f",x"26",x"87"),
  1339 => (x"d2",x"02",x"99",x"71"),
  1340 => (x"f9",x"ee",x"c1",x"87"),
  1341 => (x"f7",x"50",x"c0",x"48"),
  1342 => (x"c3",x"d3",x"c1",x"80"),
  1343 => (x"dd",x"ed",x"c1",x"40"),
  1344 => (x"c1",x"87",x"ce",x"78"),
  1345 => (x"c1",x"48",x"f5",x"ee"),
  1346 => (x"fc",x"78",x"d6",x"ed"),
  1347 => (x"e2",x"d3",x"c1",x"80"),
  1348 => (x"0e",x"4f",x"26",x"78"),
  1349 => (x"0e",x"5c",x"5b",x"5e"),
  1350 => (x"cb",x"4a",x"4c",x"71"),
  1351 => (x"e4",x"ed",x"c1",x"92"),
  1352 => (x"49",x"a2",x"c8",x"82"),
  1353 => (x"97",x"4b",x"a2",x"c9"),
  1354 => (x"97",x"1e",x"4b",x"6b"),
  1355 => (x"ca",x"1e",x"49",x"69"),
  1356 => (x"c0",x"49",x"12",x"82"),
  1357 => (x"c0",x"87",x"c6",x"e9"),
  1358 => (x"87",x"d0",x"d4",x"49"),
  1359 => (x"fb",x"c0",x"49",x"74"),
  1360 => (x"8e",x"f8",x"87",x"cd"),
  1361 => (x"1e",x"87",x"cc",x"f2"),
  1362 => (x"4b",x"71",x"1e",x"73"),
  1363 => (x"87",x"c3",x"ff",x"49"),
  1364 => (x"fe",x"fe",x"49",x"73"),
  1365 => (x"87",x"fd",x"f1",x"87"),
  1366 => (x"71",x"1e",x"73",x"1e"),
  1367 => (x"4a",x"a3",x"c6",x"4b"),
  1368 => (x"c1",x"87",x"db",x"02"),
  1369 => (x"87",x"d6",x"02",x"8a"),
  1370 => (x"da",x"c1",x"02",x"8a"),
  1371 => (x"c0",x"02",x"8a",x"87"),
  1372 => (x"02",x"8a",x"87",x"fc"),
  1373 => (x"8a",x"87",x"e1",x"c0"),
  1374 => (x"c1",x"87",x"cb",x"02"),
  1375 => (x"49",x"c7",x"87",x"db"),
  1376 => (x"c1",x"87",x"c0",x"fd"),
  1377 => (x"c7",x"c4",x"87",x"de"),
  1378 => (x"c1",x"02",x"bf",x"c0"),
  1379 => (x"c1",x"48",x"87",x"cb"),
  1380 => (x"c4",x"c7",x"c4",x"88"),
  1381 => (x"87",x"c1",x"c1",x"58"),
  1382 => (x"bf",x"c4",x"c7",x"c4"),
  1383 => (x"87",x"f9",x"c0",x"02"),
  1384 => (x"bf",x"c0",x"c7",x"c4"),
  1385 => (x"c4",x"80",x"c1",x"48"),
  1386 => (x"c0",x"58",x"c4",x"c7"),
  1387 => (x"c7",x"c4",x"87",x"eb"),
  1388 => (x"c6",x"49",x"bf",x"c0"),
  1389 => (x"c4",x"c7",x"c4",x"89"),
  1390 => (x"a9",x"b7",x"c0",x"59"),
  1391 => (x"c4",x"87",x"da",x"03"),
  1392 => (x"c0",x"48",x"c0",x"c7"),
  1393 => (x"c4",x"87",x"d2",x"78"),
  1394 => (x"02",x"bf",x"c4",x"c7"),
  1395 => (x"c7",x"c4",x"87",x"cb"),
  1396 => (x"c6",x"48",x"bf",x"c0"),
  1397 => (x"c4",x"c7",x"c4",x"80"),
  1398 => (x"d1",x"49",x"c0",x"58"),
  1399 => (x"49",x"73",x"87",x"ee"),
  1400 => (x"87",x"eb",x"f8",x"c0"),
  1401 => (x"0e",x"87",x"ee",x"ef"),
  1402 => (x"0e",x"5c",x"5b",x"5e"),
  1403 => (x"66",x"cc",x"4c",x"71"),
  1404 => (x"cb",x"4b",x"74",x"1e"),
  1405 => (x"e4",x"ed",x"c1",x"93"),
  1406 => (x"4a",x"a3",x"c4",x"83"),
  1407 => (x"eb",x"fe",x"49",x"6a"),
  1408 => (x"d2",x"c1",x"87",x"c7"),
  1409 => (x"a3",x"c8",x"7b",x"c1"),
  1410 => (x"51",x"66",x"d4",x"49"),
  1411 => (x"d8",x"49",x"a3",x"c9"),
  1412 => (x"a3",x"ca",x"51",x"66"),
  1413 => (x"51",x"66",x"dc",x"49"),
  1414 => (x"87",x"f7",x"ee",x"26"),
  1415 => (x"5c",x"5b",x"5e",x"0e"),
  1416 => (x"d0",x"ff",x"0e",x"5d"),
  1417 => (x"59",x"a6",x"d8",x"86"),
  1418 => (x"c0",x"48",x"a6",x"c4"),
  1419 => (x"c1",x"80",x"c4",x"78"),
  1420 => (x"c4",x"78",x"66",x"c4"),
  1421 => (x"c4",x"78",x"c1",x"80"),
  1422 => (x"c4",x"78",x"c1",x"80"),
  1423 => (x"c1",x"48",x"c4",x"c7"),
  1424 => (x"fc",x"c6",x"c4",x"78"),
  1425 => (x"a8",x"de",x"48",x"bf"),
  1426 => (x"f3",x"87",x"cb",x"05"),
  1427 => (x"49",x"70",x"87",x"e5"),
  1428 => (x"ce",x"59",x"a6",x"c8"),
  1429 => (x"c1",x"e6",x"87",x"fe"),
  1430 => (x"87",x"e3",x"e6",x"87"),
  1431 => (x"70",x"87",x"f0",x"e5"),
  1432 => (x"ac",x"fb",x"c0",x"4c"),
  1433 => (x"87",x"d0",x"c1",x"02"),
  1434 => (x"c1",x"05",x"66",x"d4"),
  1435 => (x"1e",x"c0",x"87",x"c2"),
  1436 => (x"c1",x"1e",x"c1",x"1e"),
  1437 => (x"c0",x"1e",x"d7",x"ef"),
  1438 => (x"87",x"eb",x"fd",x"49"),
  1439 => (x"4a",x"66",x"d0",x"c1"),
  1440 => (x"49",x"6a",x"82",x"c4"),
  1441 => (x"51",x"74",x"81",x"c7"),
  1442 => (x"1e",x"d8",x"1e",x"c1"),
  1443 => (x"81",x"c8",x"49",x"6a"),
  1444 => (x"d8",x"87",x"c0",x"e6"),
  1445 => (x"66",x"c4",x"c1",x"86"),
  1446 => (x"01",x"a8",x"c0",x"48"),
  1447 => (x"a6",x"c4",x"87",x"c7"),
  1448 => (x"ce",x"78",x"c1",x"48"),
  1449 => (x"66",x"c4",x"c1",x"87"),
  1450 => (x"cc",x"88",x"c1",x"48"),
  1451 => (x"87",x"c3",x"58",x"a6"),
  1452 => (x"cc",x"87",x"cc",x"e5"),
  1453 => (x"78",x"c2",x"48",x"a6"),
  1454 => (x"cd",x"02",x"9c",x"74"),
  1455 => (x"66",x"c4",x"87",x"d2"),
  1456 => (x"66",x"c8",x"c1",x"48"),
  1457 => (x"c7",x"cd",x"03",x"a8"),
  1458 => (x"48",x"a6",x"d8",x"87"),
  1459 => (x"fe",x"e3",x"78",x"c0"),
  1460 => (x"c1",x"4c",x"70",x"87"),
  1461 => (x"c2",x"05",x"ac",x"d0"),
  1462 => (x"66",x"d8",x"87",x"d6"),
  1463 => (x"87",x"e2",x"e6",x"7e"),
  1464 => (x"a6",x"dc",x"49",x"70"),
  1465 => (x"87",x"e7",x"e3",x"59"),
  1466 => (x"ec",x"c0",x"4c",x"70"),
  1467 => (x"ea",x"c1",x"05",x"ac"),
  1468 => (x"49",x"66",x"c4",x"87"),
  1469 => (x"c0",x"c1",x"91",x"cb"),
  1470 => (x"a1",x"c4",x"81",x"66"),
  1471 => (x"c8",x"4d",x"6a",x"4a"),
  1472 => (x"66",x"d8",x"4a",x"a1"),
  1473 => (x"c3",x"d3",x"c1",x"52"),
  1474 => (x"87",x"c3",x"e3",x"79"),
  1475 => (x"02",x"9c",x"4c",x"70"),
  1476 => (x"fb",x"c0",x"87",x"d8"),
  1477 => (x"87",x"d2",x"02",x"ac"),
  1478 => (x"f2",x"e2",x"55",x"74"),
  1479 => (x"9c",x"4c",x"70",x"87"),
  1480 => (x"c0",x"87",x"c7",x"02"),
  1481 => (x"ff",x"05",x"ac",x"fb"),
  1482 => (x"e0",x"c0",x"87",x"ee"),
  1483 => (x"55",x"c1",x"c2",x"55"),
  1484 => (x"d4",x"7d",x"97",x"c0"),
  1485 => (x"a9",x"6e",x"49",x"66"),
  1486 => (x"c4",x"87",x"db",x"05"),
  1487 => (x"66",x"c8",x"48",x"66"),
  1488 => (x"87",x"ca",x"04",x"a8"),
  1489 => (x"c1",x"48",x"66",x"c4"),
  1490 => (x"58",x"a6",x"c8",x"80"),
  1491 => (x"66",x"c8",x"87",x"c8"),
  1492 => (x"cc",x"88",x"c1",x"48"),
  1493 => (x"f6",x"e1",x"58",x"a6"),
  1494 => (x"c1",x"4c",x"70",x"87"),
  1495 => (x"c8",x"05",x"ac",x"d0"),
  1496 => (x"48",x"66",x"d0",x"87"),
  1497 => (x"a6",x"d4",x"80",x"c1"),
  1498 => (x"ac",x"d0",x"c1",x"58"),
  1499 => (x"87",x"ea",x"fd",x"02"),
  1500 => (x"d4",x"48",x"a6",x"dc"),
  1501 => (x"66",x"d8",x"78",x"66"),
  1502 => (x"a8",x"66",x"dc",x"48"),
  1503 => (x"87",x"e2",x"c9",x"05"),
  1504 => (x"48",x"a6",x"e0",x"c0"),
  1505 => (x"c4",x"78",x"f0",x"c0"),
  1506 => (x"78",x"66",x"cc",x"80"),
  1507 => (x"78",x"c0",x"80",x"c4"),
  1508 => (x"c0",x"48",x"74",x"7e"),
  1509 => (x"f0",x"c0",x"88",x"fb"),
  1510 => (x"98",x"70",x"58",x"a6"),
  1511 => (x"87",x"dd",x"c8",x"02"),
  1512 => (x"c0",x"88",x"cb",x"48"),
  1513 => (x"70",x"58",x"a6",x"f0"),
  1514 => (x"e9",x"c0",x"02",x"98"),
  1515 => (x"88",x"c9",x"48",x"87"),
  1516 => (x"58",x"a6",x"f0",x"c0"),
  1517 => (x"c3",x"02",x"98",x"70"),
  1518 => (x"c4",x"48",x"87",x"e5"),
  1519 => (x"a6",x"f0",x"c0",x"88"),
  1520 => (x"02",x"98",x"70",x"58"),
  1521 => (x"c1",x"48",x"87",x"de"),
  1522 => (x"a6",x"f0",x"c0",x"88"),
  1523 => (x"02",x"98",x"70",x"58"),
  1524 => (x"c7",x"87",x"cc",x"c3"),
  1525 => (x"e0",x"c0",x"87",x"e1"),
  1526 => (x"78",x"c0",x"48",x"a6"),
  1527 => (x"c1",x"48",x"66",x"cc"),
  1528 => (x"58",x"a6",x"d0",x"80"),
  1529 => (x"87",x"e7",x"df",x"ff"),
  1530 => (x"ec",x"c0",x"4c",x"70"),
  1531 => (x"87",x"d5",x"02",x"ac"),
  1532 => (x"02",x"66",x"e0",x"c0"),
  1533 => (x"e4",x"c0",x"87",x"c6"),
  1534 => (x"87",x"c9",x"5c",x"a6"),
  1535 => (x"f0",x"c0",x"48",x"74"),
  1536 => (x"a6",x"e8",x"c0",x"88"),
  1537 => (x"ac",x"ec",x"c0",x"58"),
  1538 => (x"ff",x"87",x"cd",x"02"),
  1539 => (x"70",x"87",x"c0",x"df"),
  1540 => (x"ac",x"ec",x"c0",x"4c"),
  1541 => (x"87",x"f3",x"ff",x"05"),
  1542 => (x"1e",x"66",x"e0",x"c0"),
  1543 => (x"1e",x"49",x"66",x"d4"),
  1544 => (x"1e",x"66",x"ec",x"c0"),
  1545 => (x"1e",x"d7",x"ef",x"c1"),
  1546 => (x"f6",x"49",x"66",x"d4"),
  1547 => (x"1e",x"c0",x"87",x"f9"),
  1548 => (x"66",x"dc",x"1e",x"ca"),
  1549 => (x"c1",x"91",x"cb",x"49"),
  1550 => (x"d8",x"81",x"66",x"d8"),
  1551 => (x"a1",x"c4",x"48",x"a6"),
  1552 => (x"bf",x"66",x"d8",x"78"),
  1553 => (x"ca",x"df",x"ff",x"49"),
  1554 => (x"c0",x"86",x"d8",x"87"),
  1555 => (x"c1",x"06",x"a8",x"b7"),
  1556 => (x"1e",x"c1",x"87",x"c8"),
  1557 => (x"66",x"c8",x"1e",x"de"),
  1558 => (x"de",x"ff",x"49",x"bf"),
  1559 => (x"86",x"c8",x"87",x"f5"),
  1560 => (x"c0",x"48",x"49",x"70"),
  1561 => (x"e4",x"c0",x"88",x"08"),
  1562 => (x"b7",x"c0",x"58",x"a6"),
  1563 => (x"e9",x"c0",x"06",x"a8"),
  1564 => (x"66",x"e0",x"c0",x"87"),
  1565 => (x"a8",x"b7",x"dd",x"48"),
  1566 => (x"6e",x"87",x"df",x"03"),
  1567 => (x"e0",x"c0",x"49",x"bf"),
  1568 => (x"e0",x"c0",x"81",x"66"),
  1569 => (x"c1",x"49",x"66",x"51"),
  1570 => (x"81",x"bf",x"6e",x"81"),
  1571 => (x"c0",x"51",x"c1",x"c2"),
  1572 => (x"c2",x"49",x"66",x"e0"),
  1573 => (x"81",x"bf",x"6e",x"81"),
  1574 => (x"7e",x"c1",x"51",x"c0"),
  1575 => (x"ff",x"87",x"de",x"c4"),
  1576 => (x"c0",x"87",x"df",x"df"),
  1577 => (x"ff",x"58",x"a6",x"e4"),
  1578 => (x"c0",x"87",x"d7",x"df"),
  1579 => (x"c0",x"58",x"a6",x"e8"),
  1580 => (x"c0",x"05",x"a8",x"ec"),
  1581 => (x"e4",x"c0",x"87",x"cb"),
  1582 => (x"e0",x"c0",x"48",x"a6"),
  1583 => (x"c4",x"c0",x"78",x"66"),
  1584 => (x"ca",x"dc",x"ff",x"87"),
  1585 => (x"49",x"66",x"c4",x"87"),
  1586 => (x"c0",x"c1",x"91",x"cb"),
  1587 => (x"80",x"71",x"48",x"66"),
  1588 => (x"4a",x"6e",x"7e",x"70"),
  1589 => (x"49",x"6e",x"82",x"c8"),
  1590 => (x"e0",x"c0",x"81",x"ca"),
  1591 => (x"e4",x"c0",x"51",x"66"),
  1592 => (x"81",x"c1",x"49",x"66"),
  1593 => (x"89",x"66",x"e0",x"c0"),
  1594 => (x"30",x"71",x"48",x"c1"),
  1595 => (x"89",x"c1",x"49",x"70"),
  1596 => (x"c4",x"7a",x"97",x"71"),
  1597 => (x"49",x"bf",x"f1",x"ca"),
  1598 => (x"29",x"66",x"e0",x"c0"),
  1599 => (x"48",x"4a",x"6a",x"97"),
  1600 => (x"f0",x"c0",x"98",x"71"),
  1601 => (x"49",x"6e",x"58",x"a6"),
  1602 => (x"4d",x"69",x"81",x"c4"),
  1603 => (x"d8",x"48",x"66",x"dc"),
  1604 => (x"c0",x"02",x"a8",x"66"),
  1605 => (x"a6",x"d8",x"87",x"c8"),
  1606 => (x"c0",x"78",x"c0",x"48"),
  1607 => (x"a6",x"d8",x"87",x"c5"),
  1608 => (x"d8",x"78",x"c1",x"48"),
  1609 => (x"e0",x"c0",x"1e",x"66"),
  1610 => (x"ff",x"49",x"75",x"1e"),
  1611 => (x"c8",x"87",x"e4",x"db"),
  1612 => (x"c0",x"4c",x"70",x"86"),
  1613 => (x"c1",x"06",x"ac",x"b7"),
  1614 => (x"85",x"74",x"87",x"d4"),
  1615 => (x"74",x"49",x"e0",x"c0"),
  1616 => (x"c1",x"4b",x"75",x"89"),
  1617 => (x"71",x"4a",x"c9",x"e9"),
  1618 => (x"87",x"ed",x"dd",x"fe"),
  1619 => (x"e8",x"c0",x"85",x"c2"),
  1620 => (x"80",x"c1",x"48",x"66"),
  1621 => (x"58",x"a6",x"ec",x"c0"),
  1622 => (x"49",x"66",x"ec",x"c0"),
  1623 => (x"a9",x"70",x"81",x"c1"),
  1624 => (x"87",x"c8",x"c0",x"02"),
  1625 => (x"c0",x"48",x"a6",x"d8"),
  1626 => (x"87",x"c5",x"c0",x"78"),
  1627 => (x"c1",x"48",x"a6",x"d8"),
  1628 => (x"1e",x"66",x"d8",x"78"),
  1629 => (x"c0",x"49",x"a4",x"c2"),
  1630 => (x"88",x"71",x"48",x"e0"),
  1631 => (x"75",x"1e",x"49",x"70"),
  1632 => (x"ce",x"da",x"ff",x"49"),
  1633 => (x"c0",x"86",x"c8",x"87"),
  1634 => (x"ff",x"01",x"a8",x"b7"),
  1635 => (x"e8",x"c0",x"87",x"c0"),
  1636 => (x"d1",x"c0",x"02",x"66"),
  1637 => (x"c9",x"49",x"6e",x"87"),
  1638 => (x"66",x"e8",x"c0",x"81"),
  1639 => (x"c1",x"48",x"6e",x"51"),
  1640 => (x"c0",x"78",x"d3",x"d4"),
  1641 => (x"49",x"6e",x"87",x"cc"),
  1642 => (x"51",x"c2",x"81",x"c9"),
  1643 => (x"d5",x"c1",x"48",x"6e"),
  1644 => (x"7e",x"c1",x"78",x"c7"),
  1645 => (x"ff",x"87",x"c6",x"c0"),
  1646 => (x"70",x"87",x"c4",x"d9"),
  1647 => (x"c0",x"02",x"6e",x"4c"),
  1648 => (x"66",x"c4",x"87",x"f5"),
  1649 => (x"a8",x"66",x"c8",x"48"),
  1650 => (x"87",x"cb",x"c0",x"04"),
  1651 => (x"c1",x"48",x"66",x"c4"),
  1652 => (x"58",x"a6",x"c8",x"80"),
  1653 => (x"c8",x"87",x"e0",x"c0"),
  1654 => (x"88",x"c1",x"48",x"66"),
  1655 => (x"c0",x"58",x"a6",x"cc"),
  1656 => (x"c6",x"c1",x"87",x"d5"),
  1657 => (x"c8",x"c0",x"05",x"ac"),
  1658 => (x"48",x"66",x"cc",x"87"),
  1659 => (x"a6",x"d0",x"80",x"c1"),
  1660 => (x"ca",x"d8",x"ff",x"58"),
  1661 => (x"d0",x"4c",x"70",x"87"),
  1662 => (x"80",x"c1",x"48",x"66"),
  1663 => (x"74",x"58",x"a6",x"d4"),
  1664 => (x"cb",x"c0",x"02",x"9c"),
  1665 => (x"48",x"66",x"c4",x"87"),
  1666 => (x"a8",x"66",x"c8",x"c1"),
  1667 => (x"87",x"f9",x"f2",x"04"),
  1668 => (x"87",x"e2",x"d7",x"ff"),
  1669 => (x"c7",x"48",x"66",x"c4"),
  1670 => (x"e5",x"c0",x"03",x"a8"),
  1671 => (x"c4",x"c7",x"c4",x"87"),
  1672 => (x"c4",x"78",x"c0",x"48"),
  1673 => (x"91",x"cb",x"49",x"66"),
  1674 => (x"81",x"66",x"c0",x"c1"),
  1675 => (x"6a",x"4a",x"a1",x"c4"),
  1676 => (x"79",x"52",x"c0",x"4a"),
  1677 => (x"c1",x"48",x"66",x"c4"),
  1678 => (x"58",x"a6",x"c8",x"80"),
  1679 => (x"ff",x"04",x"a8",x"c7"),
  1680 => (x"d0",x"ff",x"87",x"db"),
  1681 => (x"c8",x"de",x"ff",x"8e"),
  1682 => (x"00",x"20",x"3a",x"87"),
  1683 => (x"71",x"1e",x"73",x"1e"),
  1684 => (x"c6",x"02",x"9b",x"4b"),
  1685 => (x"c0",x"c7",x"c4",x"87"),
  1686 => (x"c7",x"78",x"c0",x"48"),
  1687 => (x"c0",x"c7",x"c4",x"1e"),
  1688 => (x"c1",x"1e",x"49",x"bf"),
  1689 => (x"c4",x"1e",x"e4",x"ed"),
  1690 => (x"49",x"bf",x"fc",x"c6"),
  1691 => (x"cc",x"87",x"ed",x"ee"),
  1692 => (x"fc",x"c6",x"c4",x"86"),
  1693 => (x"f2",x"e9",x"49",x"bf"),
  1694 => (x"02",x"9b",x"73",x"87"),
  1695 => (x"ed",x"c1",x"87",x"c8"),
  1696 => (x"e7",x"c0",x"49",x"e4"),
  1697 => (x"dd",x"ff",x"87",x"db"),
  1698 => (x"73",x"1e",x"87",x"cb"),
  1699 => (x"c3",x"4b",x"c0",x"1e"),
  1700 => (x"c0",x"48",x"fc",x"f7"),
  1701 => (x"c7",x"ef",x"c1",x"50"),
  1702 => (x"c8",x"c2",x"49",x"bf"),
  1703 => (x"98",x"70",x"87",x"e6"),
  1704 => (x"c1",x"87",x"c4",x"05"),
  1705 => (x"73",x"4b",x"ed",x"ea"),
  1706 => (x"e8",x"dc",x"ff",x"48"),
  1707 => (x"4d",x"4f",x"52",x"87"),
  1708 => (x"61",x"6f",x"6c",x"20"),
  1709 => (x"67",x"6e",x"69",x"64"),
  1710 => (x"69",x"61",x"66",x"20"),
  1711 => (x"00",x"64",x"65",x"6c"),
  1712 => (x"87",x"f2",x"c7",x"1e"),
  1713 => (x"c3",x"fe",x"49",x"c1"),
  1714 => (x"ed",x"e6",x"fe",x"87"),
  1715 => (x"02",x"98",x"70",x"87"),
  1716 => (x"ef",x"fe",x"87",x"cd"),
  1717 => (x"98",x"70",x"87",x"ea"),
  1718 => (x"c1",x"87",x"c4",x"02"),
  1719 => (x"c0",x"87",x"c2",x"4a"),
  1720 => (x"05",x"9a",x"72",x"4a"),
  1721 => (x"1e",x"c0",x"87",x"ce"),
  1722 => (x"49",x"d4",x"ec",x"c1"),
  1723 => (x"87",x"c1",x"f3",x"c0"),
  1724 => (x"87",x"fe",x"86",x"c4"),
  1725 => (x"87",x"ee",x"cc",x"c2"),
  1726 => (x"ec",x"c1",x"1e",x"c0"),
  1727 => (x"f2",x"c0",x"49",x"df"),
  1728 => (x"1e",x"c0",x"87",x"ef"),
  1729 => (x"70",x"87",x"c3",x"fe"),
  1730 => (x"e4",x"f2",x"c0",x"49"),
  1731 => (x"87",x"e5",x"c3",x"87"),
  1732 => (x"4f",x"26",x"8e",x"f8"),
  1733 => (x"66",x"20",x"44",x"53"),
  1734 => (x"65",x"6c",x"69",x"61"),
  1735 => (x"42",x"00",x"2e",x"64"),
  1736 => (x"69",x"74",x"6f",x"6f"),
  1737 => (x"2e",x"2e",x"67",x"6e"),
  1738 => (x"c1",x"1e",x"00",x"2e"),
  1739 => (x"c0",x"87",x"c2",x"fc"),
  1740 => (x"c1",x"87",x"cc",x"e9"),
  1741 => (x"c2",x"87",x"fa",x"fb"),
  1742 => (x"ee",x"87",x"f8",x"c0"),
  1743 => (x"1e",x"4f",x"26",x"87"),
  1744 => (x"48",x"c0",x"c7",x"c4"),
  1745 => (x"c6",x"c4",x"78",x"c0"),
  1746 => (x"78",x"c0",x"48",x"fc"),
  1747 => (x"ff",x"87",x"f1",x"fd"),
  1748 => (x"48",x"c0",x"87",x"d8"),
  1749 => (x"20",x"80",x"4f",x"26"),
  1750 => (x"74",x"69",x"78",x"45"),
  1751 => (x"42",x"20",x"80",x"00"),
  1752 => (x"00",x"6b",x"63",x"61"),
  1753 => (x"00",x"00",x"14",x"c3"),
  1754 => (x"00",x"00",x"41",x"d5"),
  1755 => (x"c3",x"00",x"00",x"00"),
  1756 => (x"f3",x"00",x"00",x"14"),
  1757 => (x"00",x"00",x"00",x"41"),
  1758 => (x"14",x"c3",x"00",x"00"),
  1759 => (x"42",x"11",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"14",x"c3",x"00"),
  1762 => (x"00",x"42",x"2f",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"14",x"c3"),
  1765 => (x"00",x"00",x"42",x"4d"),
  1766 => (x"c3",x"00",x"00",x"00"),
  1767 => (x"6b",x"00",x"00",x"14"),
  1768 => (x"00",x"00",x"00",x"42"),
  1769 => (x"14",x"c3",x"00",x"00"),
  1770 => (x"42",x"89",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"14",x"c3",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"15",x"58"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"cb",x"00",x"00",x"00"),
  1778 => (x"4e",x"00",x"00",x"1b"),
  1779 => (x"45",x"47",x"4f",x"45"),
  1780 => (x"52",x"20",x"20",x"4f"),
  1781 => (x"4c",x"00",x"4d",x"4f"),
  1782 => (x"20",x"64",x"61",x"6f"),
  1783 => (x"1e",x"00",x"2e",x"2a"),
  1784 => (x"c0",x"48",x"f0",x"fe"),
  1785 => (x"79",x"09",x"cd",x"78"),
  1786 => (x"1e",x"4f",x"26",x"09"),
  1787 => (x"bf",x"f0",x"fe",x"1e"),
  1788 => (x"26",x"26",x"48",x"7e"),
  1789 => (x"f0",x"fe",x"1e",x"4f"),
  1790 => (x"26",x"78",x"c1",x"48"),
  1791 => (x"f0",x"fe",x"1e",x"4f"),
  1792 => (x"26",x"78",x"c0",x"48"),
  1793 => (x"4a",x"71",x"1e",x"4f"),
  1794 => (x"26",x"52",x"52",x"c0"),
  1795 => (x"5b",x"5e",x"0e",x"4f"),
  1796 => (x"f4",x"0e",x"5d",x"5c"),
  1797 => (x"97",x"4d",x"71",x"86"),
  1798 => (x"a5",x"c1",x"7e",x"6d"),
  1799 => (x"48",x"6c",x"97",x"4c"),
  1800 => (x"6e",x"58",x"a6",x"c8"),
  1801 => (x"a8",x"66",x"c4",x"48"),
  1802 => (x"ff",x"87",x"c5",x"05"),
  1803 => (x"87",x"e6",x"c0",x"48"),
  1804 => (x"c2",x"87",x"ca",x"ff"),
  1805 => (x"6c",x"97",x"49",x"a5"),
  1806 => (x"4b",x"a3",x"71",x"4b"),
  1807 => (x"97",x"4b",x"6b",x"97"),
  1808 => (x"48",x"6e",x"7e",x"6c"),
  1809 => (x"a6",x"c8",x"80",x"c1"),
  1810 => (x"cc",x"98",x"c7",x"58"),
  1811 => (x"97",x"70",x"58",x"a6"),
  1812 => (x"87",x"e1",x"fe",x"7c"),
  1813 => (x"8e",x"f4",x"48",x"73"),
  1814 => (x"4c",x"26",x"4d",x"26"),
  1815 => (x"4f",x"26",x"4b",x"26"),
  1816 => (x"5c",x"5b",x"5e",x"0e"),
  1817 => (x"71",x"86",x"f4",x"0e"),
  1818 => (x"4a",x"66",x"d8",x"4c"),
  1819 => (x"c2",x"9a",x"ff",x"c3"),
  1820 => (x"6c",x"97",x"4b",x"a4"),
  1821 => (x"49",x"a1",x"73",x"49"),
  1822 => (x"6c",x"97",x"51",x"72"),
  1823 => (x"c1",x"48",x"6e",x"7e"),
  1824 => (x"58",x"a6",x"c8",x"80"),
  1825 => (x"a6",x"cc",x"98",x"c7"),
  1826 => (x"f4",x"54",x"70",x"58"),
  1827 => (x"87",x"ca",x"ff",x"8e"),
  1828 => (x"e8",x"fd",x"1e",x"1e"),
  1829 => (x"4a",x"bf",x"e0",x"87"),
  1830 => (x"c0",x"e0",x"c0",x"49"),
  1831 => (x"87",x"cb",x"02",x"99"),
  1832 => (x"ca",x"c4",x"1e",x"72"),
  1833 => (x"f7",x"fe",x"49",x"e7"),
  1834 => (x"fc",x"86",x"c4",x"87"),
  1835 => (x"7e",x"70",x"87",x"fd"),
  1836 => (x"26",x"87",x"c2",x"fd"),
  1837 => (x"c4",x"1e",x"4f",x"26"),
  1838 => (x"fd",x"49",x"e7",x"ca"),
  1839 => (x"f2",x"c1",x"87",x"c7"),
  1840 => (x"da",x"fc",x"49",x"d0"),
  1841 => (x"87",x"d5",x"c6",x"87"),
  1842 => (x"5e",x"0e",x"4f",x"26"),
  1843 => (x"0e",x"5d",x"5c",x"5b"),
  1844 => (x"bf",x"c6",x"cb",x"c4"),
  1845 => (x"de",x"f4",x"c1",x"4a"),
  1846 => (x"72",x"4c",x"49",x"bf"),
  1847 => (x"fc",x"4d",x"71",x"bc"),
  1848 => (x"4b",x"c0",x"87",x"db"),
  1849 => (x"99",x"d0",x"49",x"74"),
  1850 => (x"75",x"87",x"d5",x"02"),
  1851 => (x"71",x"99",x"d0",x"49"),
  1852 => (x"c1",x"1e",x"c0",x"1e"),
  1853 => (x"73",x"4a",x"ec",x"fb"),
  1854 => (x"c1",x"49",x"12",x"82"),
  1855 => (x"86",x"c8",x"87",x"ca"),
  1856 => (x"83",x"2d",x"2c",x"c1"),
  1857 => (x"ff",x"04",x"ab",x"c8"),
  1858 => (x"e8",x"fb",x"87",x"da"),
  1859 => (x"de",x"f4",x"c1",x"87"),
  1860 => (x"c6",x"cb",x"c4",x"48"),
  1861 => (x"4d",x"26",x"78",x"bf"),
  1862 => (x"4b",x"26",x"4c",x"26"),
  1863 => (x"00",x"00",x"4f",x"26"),
  1864 => (x"73",x"1e",x"00",x"00"),
  1865 => (x"c0",x"4b",x"71",x"1e"),
  1866 => (x"ec",x"fb",x"c1",x"4a"),
  1867 => (x"97",x"81",x"72",x"49"),
  1868 => (x"a9",x"73",x"49",x"69"),
  1869 => (x"c1",x"87",x"c4",x"05"),
  1870 => (x"c1",x"87",x"ca",x"48"),
  1871 => (x"aa",x"b7",x"c8",x"82"),
  1872 => (x"c0",x"87",x"e6",x"04"),
  1873 => (x"87",x"d2",x"ff",x"48"),
  1874 => (x"71",x"1e",x"73",x"1e"),
  1875 => (x"d1",x"ff",x"49",x"4b"),
  1876 => (x"02",x"98",x"70",x"87"),
  1877 => (x"ff",x"87",x"ec",x"c0"),
  1878 => (x"e1",x"c8",x"48",x"d0"),
  1879 => (x"48",x"d4",x"ff",x"78"),
  1880 => (x"66",x"c8",x"78",x"c5"),
  1881 => (x"c3",x"87",x"c3",x"02"),
  1882 => (x"66",x"cc",x"78",x"e0"),
  1883 => (x"ff",x"87",x"c6",x"02"),
  1884 => (x"f0",x"c3",x"48",x"d4"),
  1885 => (x"48",x"d4",x"ff",x"78"),
  1886 => (x"d0",x"ff",x"78",x"73"),
  1887 => (x"78",x"e1",x"c8",x"48"),
  1888 => (x"fe",x"78",x"e0",x"c0"),
  1889 => (x"5e",x"0e",x"87",x"d4"),
  1890 => (x"71",x"0e",x"5c",x"5b"),
  1891 => (x"e7",x"ca",x"c4",x"4c"),
  1892 => (x"87",x"f9",x"f9",x"49"),
  1893 => (x"b7",x"c0",x"4a",x"70"),
  1894 => (x"e3",x"c2",x"04",x"aa"),
  1895 => (x"aa",x"e0",x"c3",x"87"),
  1896 => (x"c1",x"87",x"c9",x"05"),
  1897 => (x"c1",x"48",x"c9",x"f9"),
  1898 => (x"87",x"d4",x"c2",x"78"),
  1899 => (x"05",x"aa",x"f0",x"c3"),
  1900 => (x"f9",x"c1",x"87",x"c9"),
  1901 => (x"78",x"c1",x"48",x"c5"),
  1902 => (x"c1",x"87",x"f5",x"c1"),
  1903 => (x"02",x"bf",x"c9",x"f9"),
  1904 => (x"4b",x"72",x"87",x"c7"),
  1905 => (x"c2",x"b3",x"c0",x"c2"),
  1906 => (x"74",x"4b",x"72",x"87"),
  1907 => (x"87",x"d1",x"05",x"9c"),
  1908 => (x"bf",x"c5",x"f9",x"c1"),
  1909 => (x"c9",x"f9",x"c1",x"1e"),
  1910 => (x"49",x"72",x"1e",x"bf"),
  1911 => (x"c8",x"87",x"e9",x"fd"),
  1912 => (x"c5",x"f9",x"c1",x"86"),
  1913 => (x"e0",x"c0",x"02",x"bf"),
  1914 => (x"c4",x"49",x"73",x"87"),
  1915 => (x"c1",x"91",x"29",x"b7"),
  1916 => (x"73",x"81",x"ec",x"fa"),
  1917 => (x"c2",x"9a",x"cf",x"4a"),
  1918 => (x"72",x"48",x"c1",x"92"),
  1919 => (x"ff",x"4a",x"70",x"30"),
  1920 => (x"69",x"48",x"72",x"ba"),
  1921 => (x"db",x"79",x"70",x"98"),
  1922 => (x"c4",x"49",x"73",x"87"),
  1923 => (x"c1",x"91",x"29",x"b7"),
  1924 => (x"73",x"81",x"ec",x"fa"),
  1925 => (x"c2",x"9a",x"cf",x"4a"),
  1926 => (x"72",x"48",x"c3",x"92"),
  1927 => (x"48",x"4a",x"70",x"30"),
  1928 => (x"79",x"70",x"b0",x"69"),
  1929 => (x"48",x"c9",x"f9",x"c1"),
  1930 => (x"f9",x"c1",x"78",x"c0"),
  1931 => (x"78",x"c0",x"48",x"c5"),
  1932 => (x"49",x"e7",x"ca",x"c4"),
  1933 => (x"70",x"87",x"d6",x"f7"),
  1934 => (x"aa",x"b7",x"c0",x"4a"),
  1935 => (x"87",x"dd",x"fd",x"03"),
  1936 => (x"d3",x"fb",x"48",x"c0"),
  1937 => (x"00",x"00",x"00",x"87"),
  1938 => (x"00",x"00",x"00",x"00"),
  1939 => (x"1e",x"73",x"1e",x"00"),
  1940 => (x"f5",x"f9",x"4b",x"71"),
  1941 => (x"fc",x"49",x"73",x"87"),
  1942 => (x"fd",x"fa",x"87",x"ec"),
  1943 => (x"4a",x"c0",x"1e",x"87"),
  1944 => (x"91",x"c4",x"49",x"72"),
  1945 => (x"81",x"ec",x"fa",x"c1"),
  1946 => (x"82",x"c1",x"79",x"c0"),
  1947 => (x"04",x"aa",x"b7",x"d0"),
  1948 => (x"4f",x"26",x"87",x"ee"),
  1949 => (x"5c",x"5b",x"5e",x"0e"),
  1950 => (x"4d",x"71",x"0e",x"5d"),
  1951 => (x"75",x"87",x"fe",x"f5"),
  1952 => (x"2a",x"b7",x"c4",x"4a"),
  1953 => (x"ec",x"fa",x"c1",x"92"),
  1954 => (x"cf",x"4c",x"75",x"82"),
  1955 => (x"6a",x"94",x"c2",x"9c"),
  1956 => (x"2b",x"74",x"4b",x"49"),
  1957 => (x"48",x"c2",x"9b",x"c3"),
  1958 => (x"4c",x"70",x"30",x"74"),
  1959 => (x"48",x"74",x"bc",x"ff"),
  1960 => (x"7a",x"70",x"98",x"71"),
  1961 => (x"73",x"87",x"ce",x"f5"),
  1962 => (x"87",x"ea",x"f9",x"48"),
  1963 => (x"00",x"00",x"00",x"00"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"00",x"00"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"00",x"00",x"00"),
  1970 => (x"00",x"00",x"00",x"00"),
  1971 => (x"00",x"00",x"00",x"00"),
  1972 => (x"00",x"00",x"00",x"00"),
  1973 => (x"00",x"00",x"00",x"00"),
  1974 => (x"00",x"00",x"00",x"00"),
  1975 => (x"00",x"00",x"00",x"00"),
  1976 => (x"00",x"00",x"00",x"00"),
  1977 => (x"00",x"00",x"00",x"00"),
  1978 => (x"00",x"00",x"00",x"00"),
  1979 => (x"25",x"26",x"1e",x"16"),
  1980 => (x"3e",x"3d",x"36",x"2e"),
  1981 => (x"48",x"d0",x"ff",x"1e"),
  1982 => (x"71",x"78",x"e1",x"c8"),
  1983 => (x"08",x"d4",x"ff",x"48"),
  1984 => (x"1e",x"4f",x"26",x"78"),
  1985 => (x"c8",x"48",x"d0",x"ff"),
  1986 => (x"48",x"71",x"78",x"e1"),
  1987 => (x"78",x"08",x"d4",x"ff"),
  1988 => (x"ff",x"48",x"66",x"c4"),
  1989 => (x"26",x"78",x"08",x"d4"),
  1990 => (x"4a",x"71",x"1e",x"4f"),
  1991 => (x"1e",x"49",x"66",x"c4"),
  1992 => (x"de",x"ff",x"49",x"72"),
  1993 => (x"48",x"d0",x"ff",x"87"),
  1994 => (x"26",x"78",x"e0",x"c0"),
  1995 => (x"71",x"1e",x"4f",x"26"),
  1996 => (x"1e",x"66",x"c4",x"4a"),
  1997 => (x"49",x"a2",x"e0",x"c1"),
  1998 => (x"c8",x"87",x"c8",x"ff"),
  1999 => (x"b7",x"c8",x"49",x"66"),
  2000 => (x"48",x"d4",x"ff",x"29"),
  2001 => (x"d0",x"ff",x"78",x"71"),
  2002 => (x"78",x"e0",x"c0",x"48"),
  2003 => (x"1e",x"4f",x"26",x"26"),
  2004 => (x"c3",x"4a",x"d4",x"ff"),
  2005 => (x"d0",x"ff",x"7a",x"ff"),
  2006 => (x"78",x"e1",x"c8",x"48"),
  2007 => (x"ca",x"c4",x"7a",x"de"),
  2008 => (x"49",x"7a",x"bf",x"f1"),
  2009 => (x"70",x"28",x"c8",x"48"),
  2010 => (x"d0",x"48",x"71",x"7a"),
  2011 => (x"71",x"7a",x"70",x"28"),
  2012 => (x"70",x"28",x"d8",x"48"),
  2013 => (x"48",x"d0",x"ff",x"7a"),
  2014 => (x"26",x"78",x"e0",x"c0"),
  2015 => (x"5b",x"5e",x"0e",x"4f"),
  2016 => (x"71",x"0e",x"5d",x"5c"),
  2017 => (x"f1",x"ca",x"c4",x"4c"),
  2018 => (x"74",x"4b",x"4d",x"bf"),
  2019 => (x"9b",x"66",x"d0",x"2b"),
  2020 => (x"66",x"d4",x"83",x"c1"),
  2021 => (x"87",x"c2",x"04",x"ab"),
  2022 => (x"4a",x"74",x"4b",x"c0"),
  2023 => (x"72",x"49",x"66",x"d0"),
  2024 => (x"75",x"b9",x"ff",x"31"),
  2025 => (x"72",x"48",x"73",x"99"),
  2026 => (x"48",x"4a",x"70",x"30"),
  2027 => (x"ca",x"c4",x"b0",x"71"),
  2028 => (x"da",x"fe",x"58",x"f5"),
  2029 => (x"26",x"4d",x"26",x"87"),
  2030 => (x"26",x"4b",x"26",x"4c"),
  2031 => (x"d0",x"ff",x"1e",x"4f"),
  2032 => (x"78",x"c9",x"c8",x"48"),
  2033 => (x"d4",x"ff",x"48",x"71"),
  2034 => (x"4f",x"26",x"78",x"08"),
  2035 => (x"49",x"4a",x"71",x"1e"),
  2036 => (x"d0",x"ff",x"87",x"eb"),
  2037 => (x"26",x"78",x"c8",x"48"),
  2038 => (x"1e",x"73",x"1e",x"4f"),
  2039 => (x"cb",x"c4",x"4b",x"71"),
  2040 => (x"c3",x"02",x"bf",x"c1"),
  2041 => (x"87",x"eb",x"c2",x"87"),
  2042 => (x"c8",x"48",x"d0",x"ff"),
  2043 => (x"49",x"73",x"78",x"c9"),
  2044 => (x"ff",x"b1",x"e0",x"c0"),
  2045 => (x"78",x"71",x"48",x"d4"),
  2046 => (x"48",x"f5",x"ca",x"c4"),
  2047 => (x"66",x"c8",x"78",x"c0"),
  2048 => (x"c3",x"87",x"c5",x"02"),
  2049 => (x"87",x"c2",x"49",x"ff"),
  2050 => (x"ca",x"c4",x"49",x"c0"),
  2051 => (x"66",x"cc",x"59",x"fd"),
  2052 => (x"c5",x"87",x"c6",x"02"),
  2053 => (x"c4",x"4a",x"d5",x"d5"),
  2054 => (x"ff",x"ff",x"cf",x"87"),
  2055 => (x"c1",x"cb",x"c4",x"4a"),
  2056 => (x"c1",x"cb",x"c4",x"5a"),
  2057 => (x"c4",x"78",x"c1",x"48"),
  2058 => (x"26",x"4d",x"26",x"87"),
  2059 => (x"26",x"4b",x"26",x"4c"),
  2060 => (x"5b",x"5e",x"0e",x"4f"),
  2061 => (x"71",x"0e",x"5d",x"5c"),
  2062 => (x"fd",x"ca",x"c4",x"4a"),
  2063 => (x"9a",x"72",x"4c",x"bf"),
  2064 => (x"49",x"87",x"cb",x"02"),
  2065 => (x"ff",x"c1",x"91",x"c8"),
  2066 => (x"83",x"71",x"4b",x"cf"),
  2067 => (x"c3",x"c2",x"87",x"c4"),
  2068 => (x"4d",x"c0",x"4b",x"cf"),
  2069 => (x"99",x"74",x"49",x"13"),
  2070 => (x"bf",x"f9",x"ca",x"c4"),
  2071 => (x"48",x"d4",x"ff",x"b9"),
  2072 => (x"b7",x"c1",x"78",x"71"),
  2073 => (x"b7",x"c8",x"85",x"2c"),
  2074 => (x"87",x"e8",x"04",x"ad"),
  2075 => (x"bf",x"f5",x"ca",x"c4"),
  2076 => (x"c4",x"80",x"c8",x"48"),
  2077 => (x"fe",x"58",x"f9",x"ca"),
  2078 => (x"73",x"1e",x"87",x"ef"),
  2079 => (x"13",x"4b",x"71",x"1e"),
  2080 => (x"cb",x"02",x"9a",x"4a"),
  2081 => (x"fe",x"49",x"72",x"87"),
  2082 => (x"4a",x"13",x"87",x"e7"),
  2083 => (x"87",x"f5",x"05",x"9a"),
  2084 => (x"1e",x"87",x"da",x"fe"),
  2085 => (x"bf",x"f5",x"ca",x"c4"),
  2086 => (x"f5",x"ca",x"c4",x"49"),
  2087 => (x"78",x"a1",x"c1",x"48"),
  2088 => (x"a9",x"b7",x"c0",x"c4"),
  2089 => (x"ff",x"87",x"db",x"03"),
  2090 => (x"ca",x"c4",x"48",x"d4"),
  2091 => (x"c4",x"78",x"bf",x"f9"),
  2092 => (x"49",x"bf",x"f5",x"ca"),
  2093 => (x"48",x"f5",x"ca",x"c4"),
  2094 => (x"c4",x"78",x"a1",x"c1"),
  2095 => (x"04",x"a9",x"b7",x"c0"),
  2096 => (x"d0",x"ff",x"87",x"e5"),
  2097 => (x"c4",x"78",x"c8",x"48"),
  2098 => (x"c0",x"48",x"c1",x"cb"),
  2099 => (x"00",x"4f",x"26",x"78"),
  2100 => (x"00",x"00",x"00",x"00"),
  2101 => (x"00",x"00",x"00",x"00"),
  2102 => (x"5f",x"5f",x"00",x"00"),
  2103 => (x"00",x"00",x"00",x"00"),
  2104 => (x"03",x"00",x"03",x"03"),
  2105 => (x"14",x"00",x"00",x"03"),
  2106 => (x"7f",x"14",x"7f",x"7f"),
  2107 => (x"00",x"00",x"14",x"7f"),
  2108 => (x"6b",x"6b",x"2e",x"24"),
  2109 => (x"4c",x"00",x"12",x"3a"),
  2110 => (x"6c",x"18",x"36",x"6a"),
  2111 => (x"30",x"00",x"32",x"56"),
  2112 => (x"77",x"59",x"4f",x"7e"),
  2113 => (x"00",x"40",x"68",x"3a"),
  2114 => (x"03",x"07",x"04",x"00"),
  2115 => (x"00",x"00",x"00",x"00"),
  2116 => (x"63",x"3e",x"1c",x"00"),
  2117 => (x"00",x"00",x"00",x"41"),
  2118 => (x"3e",x"63",x"41",x"00"),
  2119 => (x"08",x"00",x"00",x"1c"),
  2120 => (x"1c",x"1c",x"3e",x"2a"),
  2121 => (x"00",x"08",x"2a",x"3e"),
  2122 => (x"3e",x"3e",x"08",x"08"),
  2123 => (x"00",x"00",x"08",x"08"),
  2124 => (x"60",x"e0",x"80",x"00"),
  2125 => (x"00",x"00",x"00",x"00"),
  2126 => (x"08",x"08",x"08",x"08"),
  2127 => (x"00",x"00",x"08",x"08"),
  2128 => (x"60",x"60",x"00",x"00"),
  2129 => (x"40",x"00",x"00",x"00"),
  2130 => (x"0c",x"18",x"30",x"60"),
  2131 => (x"00",x"01",x"03",x"06"),
  2132 => (x"4d",x"59",x"7f",x"3e"),
  2133 => (x"00",x"00",x"3e",x"7f"),
  2134 => (x"7f",x"7f",x"06",x"04"),
  2135 => (x"00",x"00",x"00",x"00"),
  2136 => (x"59",x"71",x"63",x"42"),
  2137 => (x"00",x"00",x"46",x"4f"),
  2138 => (x"49",x"49",x"63",x"22"),
  2139 => (x"18",x"00",x"36",x"7f"),
  2140 => (x"7f",x"13",x"16",x"1c"),
  2141 => (x"00",x"00",x"10",x"7f"),
  2142 => (x"45",x"45",x"67",x"27"),
  2143 => (x"00",x"00",x"39",x"7d"),
  2144 => (x"49",x"4b",x"7e",x"3c"),
  2145 => (x"00",x"00",x"30",x"79"),
  2146 => (x"79",x"71",x"01",x"01"),
  2147 => (x"00",x"00",x"07",x"0f"),
  2148 => (x"49",x"49",x"7f",x"36"),
  2149 => (x"00",x"00",x"36",x"7f"),
  2150 => (x"69",x"49",x"4f",x"06"),
  2151 => (x"00",x"00",x"1e",x"3f"),
  2152 => (x"66",x"66",x"00",x"00"),
  2153 => (x"00",x"00",x"00",x"00"),
  2154 => (x"66",x"e6",x"80",x"00"),
  2155 => (x"00",x"00",x"00",x"00"),
  2156 => (x"14",x"14",x"08",x"08"),
  2157 => (x"00",x"00",x"22",x"22"),
  2158 => (x"14",x"14",x"14",x"14"),
  2159 => (x"00",x"00",x"14",x"14"),
  2160 => (x"14",x"14",x"22",x"22"),
  2161 => (x"00",x"00",x"08",x"08"),
  2162 => (x"59",x"51",x"03",x"02"),
  2163 => (x"3e",x"00",x"06",x"0f"),
  2164 => (x"55",x"5d",x"41",x"7f"),
  2165 => (x"00",x"00",x"1e",x"1f"),
  2166 => (x"09",x"09",x"7f",x"7e"),
  2167 => (x"00",x"00",x"7e",x"7f"),
  2168 => (x"49",x"49",x"7f",x"7f"),
  2169 => (x"00",x"00",x"36",x"7f"),
  2170 => (x"41",x"63",x"3e",x"1c"),
  2171 => (x"00",x"00",x"41",x"41"),
  2172 => (x"63",x"41",x"7f",x"7f"),
  2173 => (x"00",x"00",x"1c",x"3e"),
  2174 => (x"49",x"49",x"7f",x"7f"),
  2175 => (x"00",x"00",x"41",x"41"),
  2176 => (x"09",x"09",x"7f",x"7f"),
  2177 => (x"00",x"00",x"01",x"01"),
  2178 => (x"49",x"41",x"7f",x"3e"),
  2179 => (x"00",x"00",x"7a",x"7b"),
  2180 => (x"08",x"08",x"7f",x"7f"),
  2181 => (x"00",x"00",x"7f",x"7f"),
  2182 => (x"7f",x"7f",x"41",x"00"),
  2183 => (x"00",x"00",x"00",x"41"),
  2184 => (x"40",x"40",x"60",x"20"),
  2185 => (x"7f",x"00",x"3f",x"7f"),
  2186 => (x"36",x"1c",x"08",x"7f"),
  2187 => (x"00",x"00",x"41",x"63"),
  2188 => (x"40",x"40",x"7f",x"7f"),
  2189 => (x"7f",x"00",x"40",x"40"),
  2190 => (x"06",x"0c",x"06",x"7f"),
  2191 => (x"7f",x"00",x"7f",x"7f"),
  2192 => (x"18",x"0c",x"06",x"7f"),
  2193 => (x"00",x"00",x"7f",x"7f"),
  2194 => (x"41",x"41",x"7f",x"3e"),
  2195 => (x"00",x"00",x"3e",x"7f"),
  2196 => (x"09",x"09",x"7f",x"7f"),
  2197 => (x"3e",x"00",x"06",x"0f"),
  2198 => (x"7f",x"61",x"41",x"7f"),
  2199 => (x"00",x"00",x"40",x"7e"),
  2200 => (x"19",x"09",x"7f",x"7f"),
  2201 => (x"00",x"00",x"66",x"7f"),
  2202 => (x"59",x"4d",x"6f",x"26"),
  2203 => (x"00",x"00",x"32",x"7b"),
  2204 => (x"7f",x"7f",x"01",x"01"),
  2205 => (x"00",x"00",x"01",x"01"),
  2206 => (x"40",x"40",x"7f",x"3f"),
  2207 => (x"00",x"00",x"3f",x"7f"),
  2208 => (x"70",x"70",x"3f",x"0f"),
  2209 => (x"7f",x"00",x"0f",x"3f"),
  2210 => (x"30",x"18",x"30",x"7f"),
  2211 => (x"41",x"00",x"7f",x"7f"),
  2212 => (x"1c",x"1c",x"36",x"63"),
  2213 => (x"01",x"41",x"63",x"36"),
  2214 => (x"7c",x"7c",x"06",x"03"),
  2215 => (x"61",x"01",x"03",x"06"),
  2216 => (x"47",x"4d",x"59",x"71"),
  2217 => (x"00",x"00",x"41",x"43"),
  2218 => (x"41",x"7f",x"7f",x"00"),
  2219 => (x"01",x"00",x"00",x"41"),
  2220 => (x"18",x"0c",x"06",x"03"),
  2221 => (x"00",x"40",x"60",x"30"),
  2222 => (x"7f",x"41",x"41",x"00"),
  2223 => (x"08",x"00",x"00",x"7f"),
  2224 => (x"06",x"03",x"06",x"0c"),
  2225 => (x"80",x"00",x"08",x"0c"),
  2226 => (x"80",x"80",x"80",x"80"),
  2227 => (x"00",x"00",x"80",x"80"),
  2228 => (x"07",x"03",x"00",x"00"),
  2229 => (x"00",x"00",x"00",x"04"),
  2230 => (x"54",x"54",x"74",x"20"),
  2231 => (x"00",x"00",x"78",x"7c"),
  2232 => (x"44",x"44",x"7f",x"7f"),
  2233 => (x"00",x"00",x"38",x"7c"),
  2234 => (x"44",x"44",x"7c",x"38"),
  2235 => (x"00",x"00",x"00",x"44"),
  2236 => (x"44",x"44",x"7c",x"38"),
  2237 => (x"00",x"00",x"7f",x"7f"),
  2238 => (x"54",x"54",x"7c",x"38"),
  2239 => (x"00",x"00",x"18",x"5c"),
  2240 => (x"05",x"7f",x"7e",x"04"),
  2241 => (x"00",x"00",x"00",x"05"),
  2242 => (x"a4",x"a4",x"bc",x"18"),
  2243 => (x"00",x"00",x"7c",x"fc"),
  2244 => (x"04",x"04",x"7f",x"7f"),
  2245 => (x"00",x"00",x"78",x"7c"),
  2246 => (x"7d",x"3d",x"00",x"00"),
  2247 => (x"00",x"00",x"00",x"40"),
  2248 => (x"fd",x"80",x"80",x"80"),
  2249 => (x"00",x"00",x"00",x"7d"),
  2250 => (x"38",x"10",x"7f",x"7f"),
  2251 => (x"00",x"00",x"44",x"6c"),
  2252 => (x"7f",x"3f",x"00",x"00"),
  2253 => (x"7c",x"00",x"00",x"40"),
  2254 => (x"0c",x"18",x"0c",x"7c"),
  2255 => (x"00",x"00",x"78",x"7c"),
  2256 => (x"04",x"04",x"7c",x"7c"),
  2257 => (x"00",x"00",x"78",x"7c"),
  2258 => (x"44",x"44",x"7c",x"38"),
  2259 => (x"00",x"00",x"38",x"7c"),
  2260 => (x"24",x"24",x"fc",x"fc"),
  2261 => (x"00",x"00",x"18",x"3c"),
  2262 => (x"24",x"24",x"3c",x"18"),
  2263 => (x"00",x"00",x"fc",x"fc"),
  2264 => (x"04",x"04",x"7c",x"7c"),
  2265 => (x"00",x"00",x"08",x"0c"),
  2266 => (x"54",x"54",x"5c",x"48"),
  2267 => (x"00",x"00",x"20",x"74"),
  2268 => (x"44",x"7f",x"3f",x"04"),
  2269 => (x"00",x"00",x"00",x"44"),
  2270 => (x"40",x"40",x"7c",x"3c"),
  2271 => (x"00",x"00",x"7c",x"7c"),
  2272 => (x"60",x"60",x"3c",x"1c"),
  2273 => (x"3c",x"00",x"1c",x"3c"),
  2274 => (x"60",x"30",x"60",x"7c"),
  2275 => (x"44",x"00",x"3c",x"7c"),
  2276 => (x"38",x"10",x"38",x"6c"),
  2277 => (x"00",x"00",x"44",x"6c"),
  2278 => (x"60",x"e0",x"bc",x"1c"),
  2279 => (x"00",x"00",x"1c",x"3c"),
  2280 => (x"5c",x"74",x"64",x"44"),
  2281 => (x"00",x"00",x"44",x"4c"),
  2282 => (x"77",x"3e",x"08",x"08"),
  2283 => (x"00",x"00",x"41",x"41"),
  2284 => (x"7f",x"7f",x"00",x"00"),
  2285 => (x"00",x"00",x"00",x"00"),
  2286 => (x"3e",x"77",x"41",x"41"),
  2287 => (x"02",x"00",x"08",x"08"),
  2288 => (x"02",x"03",x"01",x"01"),
  2289 => (x"7f",x"00",x"01",x"02"),
  2290 => (x"7f",x"7f",x"7f",x"7f"),
  2291 => (x"08",x"00",x"7f",x"7f"),
  2292 => (x"3e",x"1c",x"1c",x"08"),
  2293 => (x"7f",x"7f",x"7f",x"3e"),
  2294 => (x"1c",x"3e",x"3e",x"7f"),
  2295 => (x"00",x"08",x"08",x"1c"),
  2296 => (x"7c",x"7c",x"18",x"10"),
  2297 => (x"00",x"00",x"10",x"18"),
  2298 => (x"7c",x"7c",x"30",x"10"),
  2299 => (x"10",x"00",x"10",x"30"),
  2300 => (x"78",x"60",x"60",x"30"),
  2301 => (x"42",x"00",x"06",x"1e"),
  2302 => (x"3c",x"18",x"3c",x"66"),
  2303 => (x"78",x"00",x"42",x"66"),
  2304 => (x"c6",x"c2",x"6a",x"38"),
  2305 => (x"60",x"00",x"38",x"6c"),
  2306 => (x"00",x"60",x"00",x"00"),
  2307 => (x"0e",x"00",x"60",x"00"),
  2308 => (x"5d",x"5c",x"5b",x"5e"),
  2309 => (x"4c",x"71",x"1e",x"0e"),
  2310 => (x"bf",x"d2",x"cb",x"c4"),
  2311 => (x"c0",x"4b",x"c0",x"4d"),
  2312 => (x"02",x"ab",x"74",x"1e"),
  2313 => (x"a6",x"c4",x"87",x"c7"),
  2314 => (x"c5",x"78",x"c0",x"48"),
  2315 => (x"48",x"a6",x"c4",x"87"),
  2316 => (x"66",x"c4",x"78",x"c1"),
  2317 => (x"ee",x"49",x"73",x"1e"),
  2318 => (x"86",x"c8",x"87",x"df"),
  2319 => (x"ef",x"49",x"e0",x"c0"),
  2320 => (x"a5",x"c4",x"87",x"ef"),
  2321 => (x"f0",x"49",x"6a",x"4a"),
  2322 => (x"c6",x"f1",x"87",x"f0"),
  2323 => (x"c1",x"85",x"cb",x"87"),
  2324 => (x"ab",x"b7",x"c8",x"83"),
  2325 => (x"87",x"c7",x"ff",x"04"),
  2326 => (x"26",x"4d",x"26",x"26"),
  2327 => (x"26",x"4b",x"26",x"4c"),
  2328 => (x"4a",x"71",x"1e",x"4f"),
  2329 => (x"5a",x"d6",x"cb",x"c4"),
  2330 => (x"48",x"d6",x"cb",x"c4"),
  2331 => (x"fe",x"49",x"78",x"c7"),
  2332 => (x"4f",x"26",x"87",x"dd"),
  2333 => (x"71",x"1e",x"73",x"1e"),
  2334 => (x"aa",x"b7",x"c0",x"4a"),
  2335 => (x"c2",x"87",x"d3",x"03"),
  2336 => (x"05",x"bf",x"c8",x"e0"),
  2337 => (x"4b",x"c1",x"87",x"c4"),
  2338 => (x"4b",x"c0",x"87",x"c2"),
  2339 => (x"5b",x"cc",x"e0",x"c2"),
  2340 => (x"e0",x"c2",x"87",x"c4"),
  2341 => (x"e0",x"c2",x"5a",x"cc"),
  2342 => (x"c1",x"4a",x"bf",x"c8"),
  2343 => (x"a2",x"c0",x"c1",x"9a"),
  2344 => (x"87",x"e8",x"ec",x"49"),
  2345 => (x"e0",x"c2",x"48",x"fc"),
  2346 => (x"fe",x"78",x"bf",x"c8"),
  2347 => (x"71",x"1e",x"87",x"ef"),
  2348 => (x"1e",x"66",x"c4",x"4a"),
  2349 => (x"f5",x"e9",x"49",x"72"),
  2350 => (x"4f",x"26",x"26",x"87"),
  2351 => (x"c8",x"e0",x"c2",x"1e"),
  2352 => (x"c8",x"e6",x"49",x"bf"),
  2353 => (x"ca",x"cb",x"c4",x"87"),
  2354 => (x"78",x"bf",x"e8",x"48"),
  2355 => (x"48",x"c6",x"cb",x"c4"),
  2356 => (x"c4",x"78",x"bf",x"ec"),
  2357 => (x"4a",x"bf",x"ca",x"cb"),
  2358 => (x"99",x"ff",x"cf",x"49"),
  2359 => (x"72",x"2a",x"b7",x"ca"),
  2360 => (x"c4",x"b0",x"71",x"48"),
  2361 => (x"26",x"58",x"d2",x"cb"),
  2362 => (x"5b",x"5e",x"0e",x"4f"),
  2363 => (x"71",x"0e",x"5d",x"5c"),
  2364 => (x"87",x"c8",x"ff",x"4b"),
  2365 => (x"48",x"c5",x"cb",x"c4"),
  2366 => (x"49",x"73",x"50",x"c0"),
  2367 => (x"70",x"87",x"f5",x"e5"),
  2368 => (x"9c",x"c2",x"4c",x"49"),
  2369 => (x"c1",x"49",x"ee",x"cb"),
  2370 => (x"70",x"87",x"cf",x"d7"),
  2371 => (x"cb",x"c4",x"4d",x"49"),
  2372 => (x"05",x"bf",x"97",x"c5"),
  2373 => (x"d0",x"87",x"e3",x"c1"),
  2374 => (x"cb",x"c4",x"49",x"66"),
  2375 => (x"05",x"99",x"bf",x"ce"),
  2376 => (x"66",x"d4",x"87",x"d6"),
  2377 => (x"c6",x"cb",x"c4",x"49"),
  2378 => (x"cb",x"05",x"99",x"bf"),
  2379 => (x"e5",x"49",x"73",x"87"),
  2380 => (x"98",x"70",x"87",x"c2"),
  2381 => (x"87",x"c2",x"c1",x"02"),
  2382 => (x"ff",x"fd",x"4c",x"c1"),
  2383 => (x"c1",x"49",x"75",x"87"),
  2384 => (x"70",x"87",x"e3",x"d6"),
  2385 => (x"87",x"c6",x"02",x"98"),
  2386 => (x"48",x"c5",x"cb",x"c4"),
  2387 => (x"cb",x"c4",x"50",x"c1"),
  2388 => (x"05",x"bf",x"97",x"c5"),
  2389 => (x"c4",x"87",x"e3",x"c0"),
  2390 => (x"49",x"bf",x"ce",x"cb"),
  2391 => (x"05",x"99",x"66",x"d0"),
  2392 => (x"c4",x"87",x"d5",x"ff"),
  2393 => (x"49",x"bf",x"c6",x"cb"),
  2394 => (x"05",x"99",x"66",x"d4"),
  2395 => (x"73",x"87",x"c9",x"ff"),
  2396 => (x"87",x"c0",x"e4",x"49"),
  2397 => (x"fe",x"05",x"98",x"70"),
  2398 => (x"48",x"74",x"87",x"fe"),
  2399 => (x"0e",x"87",x"da",x"fb"),
  2400 => (x"5d",x"5c",x"5b",x"5e"),
  2401 => (x"c0",x"86",x"f4",x"0e"),
  2402 => (x"bf",x"ec",x"4c",x"4d"),
  2403 => (x"48",x"a6",x"c4",x"7e"),
  2404 => (x"bf",x"d2",x"cb",x"c4"),
  2405 => (x"c0",x"1e",x"c1",x"78"),
  2406 => (x"fd",x"49",x"c7",x"1e"),
  2407 => (x"86",x"c8",x"87",x"cb"),
  2408 => (x"cd",x"02",x"98",x"70"),
  2409 => (x"fb",x"49",x"ff",x"87"),
  2410 => (x"da",x"c1",x"87",x"ca"),
  2411 => (x"87",x"c4",x"e3",x"49"),
  2412 => (x"cb",x"c4",x"4d",x"c1"),
  2413 => (x"02",x"bf",x"97",x"c5"),
  2414 => (x"e0",x"c1",x"87",x"c4"),
  2415 => (x"cb",x"c4",x"87",x"ff"),
  2416 => (x"c2",x"4b",x"bf",x"ca"),
  2417 => (x"05",x"bf",x"c8",x"e0"),
  2418 => (x"c4",x"87",x"da",x"c1"),
  2419 => (x"c0",x"c2",x"48",x"a6"),
  2420 => (x"c3",x"78",x"c0",x"c0"),
  2421 => (x"6e",x"7e",x"cf",x"f9"),
  2422 => (x"6e",x"49",x"bf",x"97"),
  2423 => (x"70",x"80",x"c1",x"48"),
  2424 => (x"cf",x"e2",x"71",x"7e"),
  2425 => (x"02",x"98",x"70",x"87"),
  2426 => (x"66",x"c4",x"87",x"c3"),
  2427 => (x"48",x"66",x"c4",x"b3"),
  2428 => (x"c8",x"28",x"b7",x"c1"),
  2429 => (x"98",x"70",x"58",x"a6"),
  2430 => (x"87",x"db",x"ff",x"05"),
  2431 => (x"e1",x"49",x"fd",x"c3"),
  2432 => (x"fa",x"c3",x"87",x"f2"),
  2433 => (x"87",x"ec",x"e1",x"49"),
  2434 => (x"ff",x"cf",x"49",x"73"),
  2435 => (x"c0",x"1e",x"71",x"99"),
  2436 => (x"87",x"da",x"fa",x"49"),
  2437 => (x"b7",x"ca",x"49",x"73"),
  2438 => (x"c1",x"1e",x"71",x"29"),
  2439 => (x"87",x"ce",x"fa",x"49"),
  2440 => (x"c7",x"c6",x"86",x"c8"),
  2441 => (x"ce",x"cb",x"c4",x"87"),
  2442 => (x"02",x"9b",x"4b",x"bf"),
  2443 => (x"e0",x"c2",x"87",x"df"),
  2444 => (x"c1",x"49",x"bf",x"c4"),
  2445 => (x"70",x"87",x"ef",x"d2"),
  2446 => (x"87",x"c4",x"05",x"98"),
  2447 => (x"87",x"d3",x"4b",x"c0"),
  2448 => (x"c1",x"49",x"e0",x"c2"),
  2449 => (x"c2",x"87",x"d3",x"d2"),
  2450 => (x"c6",x"58",x"c8",x"e0"),
  2451 => (x"c4",x"e0",x"c2",x"87"),
  2452 => (x"73",x"78",x"c0",x"48"),
  2453 => (x"05",x"99",x"c2",x"49"),
  2454 => (x"eb",x"c3",x"87",x"ce"),
  2455 => (x"87",x"d4",x"e0",x"49"),
  2456 => (x"99",x"c2",x"49",x"70"),
  2457 => (x"87",x"c2",x"c0",x"02"),
  2458 => (x"49",x"73",x"4c",x"fb"),
  2459 => (x"cf",x"05",x"99",x"c1"),
  2460 => (x"49",x"f4",x"c3",x"87"),
  2461 => (x"87",x"fc",x"df",x"ff"),
  2462 => (x"99",x"c2",x"49",x"70"),
  2463 => (x"87",x"c2",x"c0",x"02"),
  2464 => (x"49",x"73",x"4c",x"fa"),
  2465 => (x"ce",x"05",x"99",x"c8"),
  2466 => (x"49",x"f5",x"c3",x"87"),
  2467 => (x"87",x"e4",x"df",x"ff"),
  2468 => (x"99",x"c2",x"49",x"70"),
  2469 => (x"c4",x"87",x"d6",x"02"),
  2470 => (x"02",x"bf",x"d6",x"cb"),
  2471 => (x"48",x"87",x"ca",x"c0"),
  2472 => (x"cb",x"c4",x"88",x"c1"),
  2473 => (x"c2",x"c0",x"58",x"da"),
  2474 => (x"c1",x"4c",x"ff",x"87"),
  2475 => (x"c4",x"49",x"73",x"4d"),
  2476 => (x"ce",x"c0",x"05",x"99"),
  2477 => (x"49",x"f2",x"c3",x"87"),
  2478 => (x"87",x"f8",x"de",x"ff"),
  2479 => (x"99",x"c2",x"49",x"70"),
  2480 => (x"c4",x"87",x"dc",x"02"),
  2481 => (x"7e",x"bf",x"d6",x"cb"),
  2482 => (x"a8",x"b7",x"c7",x"48"),
  2483 => (x"87",x"cb",x"c0",x"03"),
  2484 => (x"80",x"c1",x"48",x"6e"),
  2485 => (x"58",x"da",x"cb",x"c4"),
  2486 => (x"fe",x"87",x"c2",x"c0"),
  2487 => (x"c3",x"4d",x"c1",x"4c"),
  2488 => (x"de",x"ff",x"49",x"fd"),
  2489 => (x"49",x"70",x"87",x"ce"),
  2490 => (x"c0",x"02",x"99",x"c2"),
  2491 => (x"cb",x"c4",x"87",x"d5"),
  2492 => (x"c0",x"02",x"bf",x"d6"),
  2493 => (x"cb",x"c4",x"87",x"c9"),
  2494 => (x"78",x"c0",x"48",x"d6"),
  2495 => (x"fd",x"87",x"c2",x"c0"),
  2496 => (x"c3",x"4d",x"c1",x"4c"),
  2497 => (x"dd",x"ff",x"49",x"fa"),
  2498 => (x"49",x"70",x"87",x"ea"),
  2499 => (x"c0",x"02",x"99",x"c2"),
  2500 => (x"cb",x"c4",x"87",x"d9"),
  2501 => (x"c7",x"48",x"bf",x"d6"),
  2502 => (x"c0",x"03",x"a8",x"b7"),
  2503 => (x"cb",x"c4",x"87",x"c9"),
  2504 => (x"78",x"c7",x"48",x"d6"),
  2505 => (x"fc",x"87",x"c2",x"c0"),
  2506 => (x"c0",x"4d",x"c1",x"4c"),
  2507 => (x"c0",x"03",x"ac",x"b7"),
  2508 => (x"66",x"c4",x"87",x"d1"),
  2509 => (x"82",x"d8",x"c1",x"4a"),
  2510 => (x"c6",x"c0",x"02",x"6a"),
  2511 => (x"74",x"4b",x"6a",x"87"),
  2512 => (x"c0",x"0f",x"73",x"49"),
  2513 => (x"1e",x"f0",x"c3",x"1e"),
  2514 => (x"f6",x"49",x"da",x"c1"),
  2515 => (x"86",x"c8",x"87",x"db"),
  2516 => (x"c0",x"02",x"98",x"70"),
  2517 => (x"a6",x"c8",x"87",x"e2"),
  2518 => (x"d6",x"cb",x"c4",x"48"),
  2519 => (x"66",x"c8",x"78",x"bf"),
  2520 => (x"c4",x"91",x"cb",x"49"),
  2521 => (x"80",x"71",x"48",x"66"),
  2522 => (x"bf",x"6e",x"7e",x"70"),
  2523 => (x"87",x"c8",x"c0",x"02"),
  2524 => (x"c8",x"4b",x"bf",x"6e"),
  2525 => (x"0f",x"73",x"49",x"66"),
  2526 => (x"c0",x"02",x"9d",x"75"),
  2527 => (x"cb",x"c4",x"87",x"c8"),
  2528 => (x"f2",x"49",x"bf",x"d6"),
  2529 => (x"e0",x"c2",x"87",x"c9"),
  2530 => (x"c0",x"02",x"bf",x"cc"),
  2531 => (x"c1",x"49",x"87",x"de"),
  2532 => (x"70",x"87",x"d3",x"cd"),
  2533 => (x"d3",x"c0",x"02",x"98"),
  2534 => (x"d6",x"cb",x"c4",x"87"),
  2535 => (x"ee",x"f1",x"49",x"bf"),
  2536 => (x"f3",x"49",x"c0",x"87"),
  2537 => (x"e0",x"c2",x"87",x"ce"),
  2538 => (x"78",x"c0",x"48",x"cc"),
  2539 => (x"e8",x"f2",x"8e",x"f4"),
  2540 => (x"5b",x"5e",x"0e",x"87"),
  2541 => (x"1e",x"0e",x"5d",x"5c"),
  2542 => (x"cb",x"c4",x"4c",x"71"),
  2543 => (x"c1",x"49",x"bf",x"d2"),
  2544 => (x"c1",x"4d",x"a1",x"cd"),
  2545 => (x"7e",x"69",x"81",x"d1"),
  2546 => (x"cf",x"02",x"9c",x"74"),
  2547 => (x"4b",x"a5",x"c4",x"87"),
  2548 => (x"cb",x"c4",x"7b",x"74"),
  2549 => (x"f2",x"49",x"bf",x"d2"),
  2550 => (x"7b",x"6e",x"87",x"c7"),
  2551 => (x"c4",x"05",x"9c",x"74"),
  2552 => (x"c2",x"4b",x"c0",x"87"),
  2553 => (x"73",x"4b",x"c1",x"87"),
  2554 => (x"87",x"c8",x"f2",x"49"),
  2555 => (x"c9",x"02",x"66",x"d4"),
  2556 => (x"cb",x"c1",x"49",x"87"),
  2557 => (x"4a",x"70",x"87",x"e4"),
  2558 => (x"4a",x"c0",x"87",x"c2"),
  2559 => (x"5a",x"d0",x"e0",x"c2"),
  2560 => (x"87",x"d5",x"f1",x"26"),
  2561 => (x"00",x"00",x"00",x"00"),
  2562 => (x"00",x"00",x"00",x"00"),
  2563 => (x"00",x"00",x"00",x"00"),
  2564 => (x"71",x"1e",x"73",x"1e"),
  2565 => (x"cb",x"c1",x"49",x"4b"),
  2566 => (x"f6",x"e8",x"fd",x"4a"),
  2567 => (x"1e",x"4a",x"70",x"87"),
  2568 => (x"fc",x"c0",x"49",x"72"),
  2569 => (x"ea",x"e8",x"fd",x"4a"),
  2570 => (x"26",x"49",x"70",x"87"),
  2571 => (x"48",x"66",x"c8",x"4a"),
  2572 => (x"49",x"72",x"50",x"71"),
  2573 => (x"fd",x"4a",x"fc",x"c0"),
  2574 => (x"71",x"87",x"d8",x"e8"),
  2575 => (x"49",x"66",x"c8",x"4a"),
  2576 => (x"51",x"72",x"81",x"c1"),
  2577 => (x"cb",x"c1",x"49",x"73"),
  2578 => (x"c6",x"e8",x"fd",x"4a"),
  2579 => (x"c8",x"4a",x"71",x"87"),
  2580 => (x"81",x"c2",x"49",x"66"),
  2581 => (x"87",x"c4",x"51",x"72"),
  2582 => (x"4c",x"26",x"4d",x"26"),
  2583 => (x"4f",x"26",x"4b",x"26"),
  2584 => (x"71",x"1e",x"73",x"1e"),
  2585 => (x"49",x"66",x"c8",x"4b"),
  2586 => (x"cc",x"91",x"cb",x"c1"),
  2587 => (x"49",x"a1",x"4a",x"66"),
  2588 => (x"c6",x"c1",x"4a",x"73"),
  2589 => (x"a1",x"72",x"92",x"d4"),
  2590 => (x"89",x"d6",x"c2",x"49"),
  2591 => (x"db",x"ff",x"48",x"71"),
  2592 => (x"5b",x"5e",x"0e",x"87"),
  2593 => (x"1e",x"0e",x"5d",x"5c"),
  2594 => (x"6b",x"97",x"4b",x"71"),
  2595 => (x"87",x"e4",x"c0",x"02"),
  2596 => (x"48",x"7e",x"6b",x"97"),
  2597 => (x"a8",x"b7",x"f0",x"c0"),
  2598 => (x"6e",x"87",x"d9",x"04"),
  2599 => (x"b7",x"f9",x"c0",x"48"),
  2600 => (x"87",x"d0",x"01",x"a8"),
  2601 => (x"49",x"6e",x"83",x"c1"),
  2602 => (x"ca",x"89",x"f0",x"c0"),
  2603 => (x"48",x"66",x"d4",x"91"),
  2604 => (x"87",x"c5",x"50",x"71"),
  2605 => (x"eb",x"c4",x"48",x"c0"),
  2606 => (x"02",x"6b",x"97",x"87"),
  2607 => (x"97",x"87",x"e9",x"c0"),
  2608 => (x"c0",x"48",x"7e",x"6b"),
  2609 => (x"04",x"a8",x"b7",x"f0"),
  2610 => (x"48",x"6e",x"87",x"de"),
  2611 => (x"a8",x"b7",x"f9",x"c0"),
  2612 => (x"c1",x"87",x"d5",x"01"),
  2613 => (x"c0",x"49",x"6e",x"83"),
  2614 => (x"66",x"d4",x"89",x"f0"),
  2615 => (x"a1",x"4a",x"bf",x"97"),
  2616 => (x"48",x"66",x"d4",x"49"),
  2617 => (x"87",x"c5",x"50",x"71"),
  2618 => (x"f7",x"c3",x"48",x"c0"),
  2619 => (x"02",x"6b",x"97",x"87"),
  2620 => (x"6b",x"97",x"87",x"cd"),
  2621 => (x"a9",x"fa",x"c0",x"49"),
  2622 => (x"c1",x"87",x"c4",x"05"),
  2623 => (x"c0",x"87",x"c5",x"83"),
  2624 => (x"87",x"e0",x"c3",x"48"),
  2625 => (x"c0",x"02",x"6b",x"97"),
  2626 => (x"6b",x"97",x"87",x"e7"),
  2627 => (x"f0",x"c0",x"48",x"7e"),
  2628 => (x"dc",x"04",x"a8",x"b7"),
  2629 => (x"c0",x"48",x"6e",x"87"),
  2630 => (x"01",x"a8",x"b7",x"f9"),
  2631 => (x"83",x"c1",x"87",x"d3"),
  2632 => (x"f0",x"c0",x"49",x"6e"),
  2633 => (x"d4",x"91",x"ca",x"89"),
  2634 => (x"84",x"c1",x"4c",x"66"),
  2635 => (x"c5",x"7c",x"97",x"71"),
  2636 => (x"c2",x"48",x"c0",x"87"),
  2637 => (x"6b",x"97",x"87",x"ee"),
  2638 => (x"87",x"e4",x"c0",x"02"),
  2639 => (x"48",x"7e",x"6b",x"97"),
  2640 => (x"a8",x"b7",x"f0",x"c0"),
  2641 => (x"6e",x"87",x"d9",x"04"),
  2642 => (x"b7",x"f9",x"c0",x"48"),
  2643 => (x"87",x"d0",x"01",x"a8"),
  2644 => (x"49",x"6e",x"83",x"c1"),
  2645 => (x"97",x"89",x"f0",x"c0"),
  2646 => (x"49",x"a1",x"4a",x"6c"),
  2647 => (x"87",x"c5",x"7c",x"97"),
  2648 => (x"ff",x"c1",x"48",x"c0"),
  2649 => (x"02",x"6b",x"97",x"87"),
  2650 => (x"6b",x"97",x"87",x"cd"),
  2651 => (x"a9",x"fa",x"c0",x"49"),
  2652 => (x"c1",x"87",x"c4",x"05"),
  2653 => (x"c0",x"87",x"c5",x"83"),
  2654 => (x"87",x"e8",x"c1",x"48"),
  2655 => (x"c0",x"02",x"6b",x"97"),
  2656 => (x"6b",x"97",x"87",x"e4"),
  2657 => (x"b7",x"f0",x"c0",x"4a"),
  2658 => (x"87",x"da",x"04",x"aa"),
  2659 => (x"aa",x"b7",x"f9",x"c0"),
  2660 => (x"c1",x"87",x"d3",x"01"),
  2661 => (x"c0",x"49",x"72",x"83"),
  2662 => (x"91",x"ca",x"89",x"f0"),
  2663 => (x"c2",x"4d",x"66",x"d4"),
  2664 => (x"7d",x"97",x"71",x"85"),
  2665 => (x"48",x"c0",x"87",x"c5"),
  2666 => (x"97",x"87",x"f9",x"c0"),
  2667 => (x"e4",x"c0",x"02",x"6b"),
  2668 => (x"7e",x"6b",x"97",x"87"),
  2669 => (x"b7",x"f0",x"c0",x"48"),
  2670 => (x"87",x"d9",x"04",x"a8"),
  2671 => (x"f9",x"c0",x"48",x"6e"),
  2672 => (x"d0",x"01",x"a8",x"b7"),
  2673 => (x"6e",x"83",x"c1",x"87"),
  2674 => (x"89",x"f0",x"c0",x"49"),
  2675 => (x"a1",x"4a",x"6d",x"97"),
  2676 => (x"c4",x"7d",x"97",x"49"),
  2677 => (x"cb",x"48",x"c0",x"87"),
  2678 => (x"02",x"6b",x"97",x"87"),
  2679 => (x"48",x"c0",x"87",x"c4"),
  2680 => (x"48",x"c1",x"87",x"c2"),
  2681 => (x"87",x"f0",x"f9",x"26"),
  2682 => (x"5c",x"5b",x"5e",x"0e"),
  2683 => (x"86",x"f8",x"0e",x"5d"),
  2684 => (x"4c",x"c0",x"4d",x"71"),
  2685 => (x"d2",x"cc",x"c4",x"4b"),
  2686 => (x"ee",x"cb",x"fe",x"49"),
  2687 => (x"c0",x"4a",x"70",x"87"),
  2688 => (x"c2",x"04",x"aa",x"b7"),
  2689 => (x"aa",x"ca",x"87",x"f2"),
  2690 => (x"87",x"ec",x"c2",x"02"),
  2691 => (x"02",x"aa",x"e0",x"c0"),
  2692 => (x"aa",x"c9",x"87",x"cf"),
  2693 => (x"cd",x"87",x"ca",x"02"),
  2694 => (x"87",x"c5",x"02",x"aa"),
  2695 => (x"c6",x"05",x"aa",x"ca"),
  2696 => (x"02",x"9c",x"74",x"87"),
  2697 => (x"c0",x"87",x"d1",x"c2"),
  2698 => (x"cc",x"05",x"aa",x"e2"),
  2699 => (x"c1",x"49",x"74",x"87"),
  2700 => (x"c3",x"4c",x"71",x"b9"),
  2701 => (x"fc",x"fe",x"9c",x"ff"),
  2702 => (x"05",x"9c",x"74",x"87"),
  2703 => (x"c1",x"87",x"e7",x"c1"),
  2704 => (x"04",x"aa",x"b7",x"e1"),
  2705 => (x"fa",x"c1",x"87",x"c8"),
  2706 => (x"c1",x"06",x"aa",x"b7"),
  2707 => (x"c1",x"c1",x"87",x"d8"),
  2708 => (x"c8",x"04",x"aa",x"b7"),
  2709 => (x"b7",x"da",x"c1",x"87"),
  2710 => (x"c9",x"c1",x"06",x"aa"),
  2711 => (x"b7",x"f0",x"c0",x"87"),
  2712 => (x"87",x"c8",x"04",x"aa"),
  2713 => (x"aa",x"b7",x"f9",x"c0"),
  2714 => (x"87",x"fa",x"c0",x"06"),
  2715 => (x"02",x"aa",x"db",x"c1"),
  2716 => (x"c1",x"87",x"f3",x"c0"),
  2717 => (x"c0",x"02",x"aa",x"dd"),
  2718 => (x"ed",x"c0",x"87",x"ec"),
  2719 => (x"e5",x"c0",x"02",x"aa"),
  2720 => (x"aa",x"df",x"c1",x"87"),
  2721 => (x"c0",x"87",x"df",x"02"),
  2722 => (x"d9",x"02",x"aa",x"ec"),
  2723 => (x"aa",x"fd",x"c0",x"87"),
  2724 => (x"c1",x"87",x"d3",x"02"),
  2725 => (x"cd",x"02",x"aa",x"fe"),
  2726 => (x"aa",x"fa",x"c0",x"87"),
  2727 => (x"c0",x"87",x"c7",x"02"),
  2728 => (x"fd",x"05",x"aa",x"ef"),
  2729 => (x"ff",x"c0",x"87",x"cf"),
  2730 => (x"fd",x"03",x"ab",x"b7"),
  2731 => (x"a3",x"75",x"87",x"c7"),
  2732 => (x"72",x"83",x"c1",x"49"),
  2733 => (x"87",x"fd",x"fc",x"51"),
  2734 => (x"c0",x"49",x"a3",x"75"),
  2735 => (x"03",x"aa",x"b7",x"51"),
  2736 => (x"7e",x"c4",x"87",x"c4"),
  2737 => (x"9b",x"73",x"87",x"df"),
  2738 => (x"c4",x"87",x"c7",x"05"),
  2739 => (x"78",x"c3",x"48",x"a6"),
  2740 => (x"9c",x"74",x"87",x"d0"),
  2741 => (x"c1",x"87",x"c4",x"02"),
  2742 => (x"c0",x"87",x"c2",x"7e"),
  2743 => (x"48",x"a6",x"c4",x"7e"),
  2744 => (x"66",x"c4",x"78",x"6e"),
  2745 => (x"f8",x"48",x"6e",x"7e"),
  2746 => (x"87",x"ec",x"f5",x"8e"),
  2747 => (x"5c",x"5b",x"5e",x"0e"),
  2748 => (x"4d",x"71",x"0e",x"5d"),
  2749 => (x"4b",x"da",x"cb",x"c4"),
  2750 => (x"f8",x"c0",x"4a",x"c0"),
  2751 => (x"d5",x"d7",x"fd",x"49"),
  2752 => (x"c4",x"1e",x"75",x"87"),
  2753 => (x"fd",x"49",x"d2",x"cc"),
  2754 => (x"c4",x"87",x"c3",x"fc"),
  2755 => (x"05",x"98",x"70",x"86"),
  2756 => (x"4c",x"c1",x"87",x"c5"),
  2757 => (x"c1",x"87",x"ea",x"c0"),
  2758 => (x"87",x"ea",x"c0",x"49"),
  2759 => (x"05",x"9c",x"4c",x"70"),
  2760 => (x"cb",x"c4",x"87",x"c9"),
  2761 => (x"dd",x"49",x"bf",x"de"),
  2762 => (x"74",x"4c",x"70",x"87"),
  2763 => (x"87",x"cb",x"05",x"9c"),
  2764 => (x"48",x"da",x"cb",x"c4"),
  2765 => (x"bf",x"ee",x"cb",x"c4"),
  2766 => (x"c4",x"87",x"c6",x"78"),
  2767 => (x"c0",x"48",x"de",x"cb"),
  2768 => (x"f4",x"48",x"74",x"78"),
  2769 => (x"5e",x"0e",x"87",x"d2"),
  2770 => (x"0e",x"5d",x"5c",x"5b"),
  2771 => (x"71",x"86",x"d4",x"ff"),
  2772 => (x"7e",x"97",x"c0",x"4c"),
  2773 => (x"c0",x"48",x"a6",x"c4"),
  2774 => (x"50",x"80",x"c0",x"50"),
  2775 => (x"c0",x"50",x"80",x"c0"),
  2776 => (x"c0",x"4d",x"50",x"80"),
  2777 => (x"80",x"c4",x"78",x"80"),
  2778 => (x"80",x"c4",x"78",x"c0"),
  2779 => (x"80",x"c4",x"78",x"c0"),
  2780 => (x"cc",x"c4",x"78",x"c0"),
  2781 => (x"c5",x"05",x"bf",x"da"),
  2782 => (x"d0",x"48",x"c1",x"87"),
  2783 => (x"cc",x"c4",x"87",x"c3"),
  2784 => (x"78",x"c0",x"48",x"d2"),
  2785 => (x"78",x"c0",x"80",x"d0"),
  2786 => (x"cc",x"c4",x"80",x"f4"),
  2787 => (x"c3",x"78",x"bf",x"de"),
  2788 => (x"c0",x"48",x"f3",x"c0"),
  2789 => (x"ee",x"cb",x"c4",x"78"),
  2790 => (x"c2",x"78",x"c0",x"48"),
  2791 => (x"f9",x"49",x"f3",x"ff"),
  2792 => (x"a6",x"dc",x"87",x"c6"),
  2793 => (x"02",x"a8",x"c3",x"58"),
  2794 => (x"97",x"87",x"d0",x"cd"),
  2795 => (x"02",x"9b",x"4b",x"6e"),
  2796 => (x"8b",x"c1",x"87",x"d8"),
  2797 => (x"87",x"f5",x"c1",x"02"),
  2798 => (x"e4",x"c3",x"02",x"8b"),
  2799 => (x"c7",x"02",x"8b",x"87"),
  2800 => (x"02",x"8b",x"87",x"c4"),
  2801 => (x"cc",x"87",x"c3",x"c8"),
  2802 => (x"a6",x"c4",x"87",x"f1"),
  2803 => (x"c2",x"50",x"c0",x"48"),
  2804 => (x"c2",x"4a",x"f3",x"ff"),
  2805 => (x"fd",x"49",x"e3",x"fe"),
  2806 => (x"70",x"87",x"f4",x"d1"),
  2807 => (x"87",x"c6",x"05",x"98"),
  2808 => (x"cc",x"7e",x"97",x"c1"),
  2809 => (x"ff",x"c2",x"87",x"d5"),
  2810 => (x"fe",x"c2",x"4a",x"f3"),
  2811 => (x"d1",x"fd",x"49",x"e8"),
  2812 => (x"98",x"70",x"87",x"dd"),
  2813 => (x"c2",x"87",x"c6",x"05"),
  2814 => (x"fe",x"cb",x"7e",x"97"),
  2815 => (x"f3",x"ff",x"c2",x"87"),
  2816 => (x"ee",x"fe",x"c2",x"4a"),
  2817 => (x"c6",x"d1",x"fd",x"49"),
  2818 => (x"05",x"98",x"70",x"87"),
  2819 => (x"c3",x"87",x"c6",x"c0"),
  2820 => (x"e6",x"cb",x"7e",x"97"),
  2821 => (x"f3",x"ff",x"c2",x"87"),
  2822 => (x"f5",x"fe",x"c2",x"4a"),
  2823 => (x"ee",x"d0",x"fd",x"49"),
  2824 => (x"05",x"98",x"70",x"87"),
  2825 => (x"c4",x"87",x"d4",x"cb"),
  2826 => (x"ce",x"cb",x"7e",x"97"),
  2827 => (x"66",x"97",x"c4",x"87"),
  2828 => (x"a6",x"e0",x"c0",x"48"),
  2829 => (x"05",x"98",x"70",x"58"),
  2830 => (x"c8",x"87",x"cd",x"c1"),
  2831 => (x"78",x"c0",x"48",x"a6"),
  2832 => (x"05",x"66",x"97",x"c7"),
  2833 => (x"c4",x"87",x"cd",x"c1"),
  2834 => (x"02",x"bf",x"c6",x"cc"),
  2835 => (x"ff",x"87",x"c7",x"c0"),
  2836 => (x"c0",x"50",x"c1",x"80"),
  2837 => (x"ff",x"c2",x"87",x"fe"),
  2838 => (x"cb",x"c4",x"1e",x"f3"),
  2839 => (x"f6",x"fd",x"49",x"fe"),
  2840 => (x"86",x"c4",x"87",x"ec"),
  2841 => (x"c0",x"02",x"98",x"70"),
  2842 => (x"a6",x"c7",x"87",x"c8"),
  2843 => (x"c0",x"50",x"c1",x"48"),
  2844 => (x"a6",x"c5",x"87",x"c5"),
  2845 => (x"c3",x"50",x"c4",x"48"),
  2846 => (x"c4",x"1e",x"ca",x"fa"),
  2847 => (x"fd",x"49",x"d2",x"cc"),
  2848 => (x"c4",x"87",x"e7",x"f9"),
  2849 => (x"87",x"cc",x"c0",x"86"),
  2850 => (x"c1",x"48",x"66",x"dc"),
  2851 => (x"c3",x"c0",x"05",x"a8"),
  2852 => (x"7e",x"97",x"c0",x"87"),
  2853 => (x"48",x"66",x"97",x"c4"),
  2854 => (x"a6",x"c4",x"80",x"c1"),
  2855 => (x"da",x"c9",x"50",x"08"),
  2856 => (x"48",x"a6",x"d4",x"87"),
  2857 => (x"78",x"66",x"e0",x"c0"),
  2858 => (x"48",x"66",x"97",x"c4"),
  2859 => (x"58",x"a6",x"e0",x"c0"),
  2860 => (x"c0",x"05",x"98",x"70"),
  2861 => (x"1e",x"ca",x"87",x"fb"),
  2862 => (x"ff",x"c2",x"1e",x"c0"),
  2863 => (x"d3",x"fd",x"49",x"f3"),
  2864 => (x"86",x"c8",x"87",x"cf"),
  2865 => (x"e0",x"c0",x"49",x"70"),
  2866 => (x"66",x"dc",x"59",x"a6"),
  2867 => (x"87",x"d3",x"c0",x"02"),
  2868 => (x"b7",x"e3",x"c1",x"48"),
  2869 => (x"ca",x"c0",x"01",x"a8"),
  2870 => (x"49",x"a5",x"c1",x"87"),
  2871 => (x"02",x"a9",x"66",x"dc"),
  2872 => (x"c5",x"87",x"c8",x"c0"),
  2873 => (x"50",x"c2",x"48",x"a6"),
  2874 => (x"dc",x"87",x"ce",x"c2"),
  2875 => (x"c8",x"c2",x"4d",x"66"),
  2876 => (x"48",x"66",x"dc",x"87"),
  2877 => (x"c1",x"05",x"a8",x"c1"),
  2878 => (x"ff",x"c2",x"87",x"ff"),
  2879 => (x"fe",x"c2",x"4a",x"f3"),
  2880 => (x"cd",x"fd",x"49",x"c7"),
  2881 => (x"98",x"70",x"87",x"c9"),
  2882 => (x"87",x"cf",x"c0",x"05"),
  2883 => (x"48",x"a6",x"e0",x"c0"),
  2884 => (x"78",x"f0",x"e4",x"c0"),
  2885 => (x"78",x"c0",x"80",x"c4"),
  2886 => (x"c2",x"87",x"c7",x"c1"),
  2887 => (x"c2",x"4a",x"f3",x"ff"),
  2888 => (x"fd",x"49",x"cd",x"fe"),
  2889 => (x"70",x"87",x"e8",x"cc"),
  2890 => (x"cf",x"c0",x"05",x"98"),
  2891 => (x"a6",x"e0",x"c0",x"87"),
  2892 => (x"f0",x"e4",x"c0",x"48"),
  2893 => (x"c1",x"80",x"c4",x"78"),
  2894 => (x"87",x"e6",x"c0",x"78"),
  2895 => (x"4a",x"f3",x"ff",x"c2"),
  2896 => (x"49",x"d8",x"fe",x"c2"),
  2897 => (x"87",x"c7",x"cc",x"fd"),
  2898 => (x"c0",x"05",x"98",x"70"),
  2899 => (x"e0",x"c0",x"87",x"cf"),
  2900 => (x"e0",x"c0",x"48",x"a6"),
  2901 => (x"80",x"c4",x"78",x"c0"),
  2902 => (x"c5",x"c0",x"78",x"c1"),
  2903 => (x"48",x"a6",x"c5",x"87"),
  2904 => (x"ac",x"75",x"50",x"c2"),
  2905 => (x"87",x"ce",x"c0",x"05"),
  2906 => (x"48",x"f6",x"cb",x"c4"),
  2907 => (x"78",x"66",x"e0",x"c0"),
  2908 => (x"e4",x"c0",x"80",x"fc"),
  2909 => (x"97",x"c0",x"78",x"66"),
  2910 => (x"66",x"97",x"c4",x"7e"),
  2911 => (x"c4",x"80",x"c1",x"48"),
  2912 => (x"c5",x"50",x"08",x"a6"),
  2913 => (x"e8",x"c0",x"87",x"f5"),
  2914 => (x"ff",x"c2",x"1e",x"a6"),
  2915 => (x"f0",x"eb",x"49",x"f3"),
  2916 => (x"70",x"86",x"c4",x"87"),
  2917 => (x"c8",x"c0",x"05",x"98"),
  2918 => (x"48",x"a6",x"c5",x"87"),
  2919 => (x"e3",x"c0",x"50",x"c2"),
  2920 => (x"97",x"ea",x"c0",x"87"),
  2921 => (x"c0",x"1e",x"49",x"66"),
  2922 => (x"49",x"66",x"97",x"ed"),
  2923 => (x"97",x"f0",x"c0",x"1e"),
  2924 => (x"eb",x"ea",x"49",x"66"),
  2925 => (x"70",x"86",x"c8",x"87"),
  2926 => (x"81",x"d6",x"c2",x"49"),
  2927 => (x"66",x"c8",x"48",x"71"),
  2928 => (x"58",x"a6",x"cc",x"80"),
  2929 => (x"c4",x"7e",x"97",x"c0"),
  2930 => (x"97",x"c4",x"87",x"f1"),
  2931 => (x"e0",x"c0",x"48",x"66"),
  2932 => (x"98",x"70",x"58",x"a6"),
  2933 => (x"87",x"d7",x"c0",x"05"),
  2934 => (x"1e",x"c0",x"1e",x"ca"),
  2935 => (x"49",x"f3",x"ff",x"c2"),
  2936 => (x"87",x"ed",x"ce",x"fd"),
  2937 => (x"49",x"70",x"86",x"c8"),
  2938 => (x"59",x"97",x"a6",x"ca"),
  2939 => (x"dc",x"87",x"c2",x"c4"),
  2940 => (x"a8",x"c1",x"48",x"66"),
  2941 => (x"87",x"f9",x"c3",x"05"),
  2942 => (x"1e",x"a6",x"e8",x"c0"),
  2943 => (x"49",x"f3",x"ff",x"c2"),
  2944 => (x"c4",x"87",x"fe",x"e9"),
  2945 => (x"05",x"98",x"70",x"86"),
  2946 => (x"c5",x"87",x"c8",x"c0"),
  2947 => (x"50",x"c2",x"48",x"a6"),
  2948 => (x"c0",x"87",x"db",x"c3"),
  2949 => (x"49",x"66",x"97",x"ea"),
  2950 => (x"97",x"ed",x"c0",x"1e"),
  2951 => (x"c0",x"1e",x"49",x"66"),
  2952 => (x"49",x"66",x"97",x"f0"),
  2953 => (x"c8",x"87",x"f9",x"e8"),
  2954 => (x"c6",x"7e",x"70",x"86"),
  2955 => (x"c0",x"48",x"66",x"97"),
  2956 => (x"70",x"58",x"a6",x"e0"),
  2957 => (x"e1",x"c0",x"05",x"98"),
  2958 => (x"49",x"a4",x"c1",x"87"),
  2959 => (x"ed",x"c2",x"05",x"ad"),
  2960 => (x"ee",x"cb",x"c4",x"87"),
  2961 => (x"e5",x"c2",x"05",x"bf"),
  2962 => (x"c2",x"49",x"6e",x"87"),
  2963 => (x"48",x"71",x"81",x"d6"),
  2964 => (x"c4",x"80",x"66",x"c8"),
  2965 => (x"c2",x"58",x"f2",x"cb"),
  2966 => (x"66",x"dc",x"87",x"d4"),
  2967 => (x"05",x"a8",x"c1",x"48"),
  2968 => (x"74",x"87",x"cb",x"c2"),
  2969 => (x"ce",x"c0",x"05",x"ad"),
  2970 => (x"c2",x"49",x"6e",x"87"),
  2971 => (x"48",x"71",x"81",x"d6"),
  2972 => (x"c4",x"80",x"66",x"c8"),
  2973 => (x"c1",x"58",x"ee",x"cb"),
  2974 => (x"c1",x"06",x"ad",x"b7"),
  2975 => (x"48",x"6e",x"87",x"ce"),
  2976 => (x"c0",x"88",x"66",x"cc"),
  2977 => (x"74",x"58",x"a6",x"e0"),
  2978 => (x"ce",x"c0",x"05",x"ad"),
  2979 => (x"d4",x"49",x"70",x"87"),
  2980 => (x"48",x"71",x"91",x"66"),
  2981 => (x"c4",x"80",x"66",x"d0"),
  2982 => (x"c1",x"58",x"ea",x"cb"),
  2983 => (x"05",x"ad",x"49",x"a4"),
  2984 => (x"c4",x"87",x"d8",x"c0"),
  2985 => (x"05",x"bf",x"ee",x"cb"),
  2986 => (x"6e",x"87",x"d0",x"c0"),
  2987 => (x"81",x"d6",x"c2",x"49"),
  2988 => (x"71",x"81",x"66",x"c8"),
  2989 => (x"c4",x"88",x"c1",x"48"),
  2990 => (x"dc",x"58",x"f2",x"cb"),
  2991 => (x"66",x"d4",x"49",x"66"),
  2992 => (x"d0",x"48",x"71",x"91"),
  2993 => (x"a6",x"d4",x"80",x"66"),
  2994 => (x"87",x"dd",x"c0",x"58"),
  2995 => (x"d6",x"c2",x"49",x"6e"),
  2996 => (x"91",x"66",x"d4",x"81"),
  2997 => (x"66",x"d0",x"48",x"71"),
  2998 => (x"58",x"a6",x"d4",x"80"),
  2999 => (x"c0",x"05",x"ac",x"c1"),
  3000 => (x"cb",x"c4",x"87",x"c7"),
  3001 => (x"66",x"d0",x"48",x"e6"),
  3002 => (x"48",x"a6",x"cc",x"78"),
  3003 => (x"97",x"c0",x"78",x"6e"),
  3004 => (x"66",x"97",x"c4",x"7e"),
  3005 => (x"c4",x"80",x"c1",x"48"),
  3006 => (x"d8",x"50",x"08",x"a6"),
  3007 => (x"a8",x"c4",x"48",x"66"),
  3008 => (x"87",x"c7",x"c0",x"02"),
  3009 => (x"02",x"66",x"97",x"c5"),
  3010 => (x"c7",x"87",x"d0",x"f2"),
  3011 => (x"c0",x"05",x"66",x"97"),
  3012 => (x"a6",x"c5",x"87",x"c8"),
  3013 => (x"c0",x"50",x"c4",x"48"),
  3014 => (x"ad",x"74",x"87",x"f1"),
  3015 => (x"87",x"eb",x"c0",x"05"),
  3016 => (x"bf",x"e6",x"cb",x"c4"),
  3017 => (x"c6",x"cc",x"c4",x"4a"),
  3018 => (x"88",x"72",x"48",x"bf"),
  3019 => (x"cb",x"c4",x"4a",x"70"),
  3020 => (x"72",x"49",x"bf",x"f6"),
  3021 => (x"4a",x"09",x"72",x"1e"),
  3022 => (x"87",x"e3",x"cb",x"fd"),
  3023 => (x"4a",x"26",x"49",x"70"),
  3024 => (x"bf",x"ea",x"cb",x"c4"),
  3025 => (x"c4",x"80",x"71",x"48"),
  3026 => (x"74",x"58",x"f2",x"cb"),
  3027 => (x"c0",x"03",x"ad",x"b7"),
  3028 => (x"a6",x"c5",x"87",x"c5"),
  3029 => (x"c5",x"50",x"c4",x"48"),
  3030 => (x"c0",x"02",x"66",x"97"),
  3031 => (x"cb",x"c4",x"87",x"c9"),
  3032 => (x"78",x"c0",x"48",x"de"),
  3033 => (x"c4",x"87",x"c4",x"c0"),
  3034 => (x"c0",x"5d",x"e2",x"cb"),
  3035 => (x"c4",x"1e",x"a6",x"e8"),
  3036 => (x"49",x"bf",x"ea",x"cb"),
  3037 => (x"c4",x"87",x"d9",x"e2"),
  3038 => (x"fe",x"cb",x"c4",x"86"),
  3039 => (x"66",x"97",x"c5",x"5c"),
  3040 => (x"8e",x"d4",x"ff",x"48"),
  3041 => (x"41",x"87",x"d1",x"e3"),
  3042 => (x"4f",x"49",x"44",x"55"),
  3043 => (x"44",x"4f",x"4d",x"00"),
  3044 => (x"32",x"2f",x"31",x"45"),
  3045 => (x"00",x"32",x"35",x"33"),
  3046 => (x"45",x"44",x"4f",x"4d"),
  3047 => (x"30",x"32",x"2f",x"31"),
  3048 => (x"46",x"00",x"38",x"34"),
  3049 => (x"00",x"45",x"4c",x"49"),
  3050 => (x"43",x"41",x"52",x"54"),
  3051 => (x"52",x"50",x"00",x"4b"),
  3052 => (x"50",x"41",x"47",x"45"),
  3053 => (x"44",x"4e",x"49",x"00"),
  3054 => (x"0e",x"00",x"58",x"45"),
  3055 => (x"0e",x"5c",x"5b",x"5e"),
  3056 => (x"4c",x"c1",x"4b",x"71"),
  3057 => (x"bf",x"ea",x"cb",x"c4"),
  3058 => (x"d0",x"04",x"ab",x"b7"),
  3059 => (x"ee",x"cb",x"c4",x"87"),
  3060 => (x"01",x"ab",x"b7",x"bf"),
  3061 => (x"cb",x"c4",x"87",x"c7"),
  3062 => (x"d3",x"48",x"bf",x"fa"),
  3063 => (x"ed",x"49",x"74",x"87"),
  3064 => (x"84",x"c1",x"87",x"e4"),
  3065 => (x"bf",x"de",x"cb",x"c4"),
  3066 => (x"ff",x"06",x"ac",x"b7"),
  3067 => (x"48",x"ff",x"87",x"d6"),
  3068 => (x"00",x"87",x"e7",x"e1"),
  3069 => (x"00",x"00",x"00",x"00"),
  3070 => (x"00",x"00",x"00",x"00"),
  3071 => (x"00",x"00",x"00",x"00"),
  3072 => (x"00",x"00",x"00",x"00"),
  3073 => (x"00",x"00",x"00",x"00"),
  3074 => (x"00",x"00",x"00",x"00"),
  3075 => (x"00",x"00",x"00",x"00"),
  3076 => (x"00",x"00",x"00",x"00"),
  3077 => (x"00",x"00",x"00",x"00"),
  3078 => (x"00",x"00",x"00",x"00"),
  3079 => (x"00",x"00",x"00",x"00"),
  3080 => (x"00",x"00",x"00",x"00"),
  3081 => (x"00",x"00",x"00",x"00"),
  3082 => (x"00",x"00",x"00",x"00"),
  3083 => (x"00",x"00",x"00",x"00"),
  3084 => (x"00",x"00",x"00",x"00"),
  3085 => (x"1e",x"00",x"00",x"00"),
  3086 => (x"4b",x"71",x"1e",x"73"),
  3087 => (x"49",x"72",x"1e",x"4a"),
  3088 => (x"c8",x"fd",x"4a",x"ca"),
  3089 => (x"49",x"70",x"87",x"cd"),
  3090 => (x"91",x"d0",x"4a",x"26"),
  3091 => (x"49",x"72",x"1e",x"71"),
  3092 => (x"c7",x"fd",x"4a",x"ca"),
  3093 => (x"4a",x"71",x"87",x"fd"),
  3094 => (x"a1",x"72",x"49",x"26"),
  3095 => (x"99",x"ff",x"c3",x"49"),
  3096 => (x"87",x"c4",x"48",x"71"),
  3097 => (x"4c",x"26",x"4d",x"26"),
  3098 => (x"4f",x"26",x"4b",x"26"),
  3099 => (x"71",x"1e",x"73",x"1e"),
  3100 => (x"c4",x"49",x"4a",x"4b"),
  3101 => (x"91",x"ca",x"29",x"b7"),
  3102 => (x"a1",x"72",x"9a",x"cf"),
  3103 => (x"99",x"ff",x"c3",x"49"),
  3104 => (x"87",x"e4",x"48",x"71"),
  3105 => (x"71",x"1e",x"73",x"1e"),
  3106 => (x"87",x"e0",x"49",x"4a"),
  3107 => (x"9b",x"4b",x"49",x"70"),
  3108 => (x"c1",x"87",x"c2",x"05"),
  3109 => (x"de",x"cb",x"c4",x"4b"),
  3110 => (x"06",x"ab",x"b7",x"bf"),
  3111 => (x"73",x"4b",x"87",x"c1"),
  3112 => (x"87",x"e2",x"ea",x"49"),
  3113 => (x"ff",x"fe",x"48",x"73"),
  3114 => (x"f1",x"c4",x"1e",x"87"),
  3115 => (x"c4",x"59",x"97",x"da"),
  3116 => (x"c4",x"48",x"d7",x"f1"),
  3117 => (x"66",x"c8",x"50",x"66"),
  3118 => (x"50",x"66",x"cc",x"50"),
  3119 => (x"73",x"1e",x"4f",x"26"),
  3120 => (x"ff",x"4b",x"71",x"1e"),
  3121 => (x"c5",x"c8",x"48",x"d0"),
  3122 => (x"48",x"d4",x"ff",x"78"),
  3123 => (x"73",x"78",x"e1",x"c1"),
  3124 => (x"b7",x"c8",x"4a",x"49"),
  3125 => (x"c3",x"78",x"72",x"2a"),
  3126 => (x"78",x"71",x"99",x"ff"),
  3127 => (x"c4",x"48",x"d0",x"ff"),
  3128 => (x"87",x"c4",x"fe",x"78"),
  3129 => (x"d4",x"f2",x"c4",x"1e"),
  3130 => (x"f1",x"c4",x"59",x"9f"),
  3131 => (x"78",x"c1",x"48",x"e4"),
  3132 => (x"5e",x"0e",x"4f",x"26"),
  3133 => (x"71",x"0e",x"5c",x"5b"),
  3134 => (x"48",x"d0",x"ff",x"4c"),
  3135 => (x"ff",x"78",x"c5",x"c8"),
  3136 => (x"e4",x"c1",x"48",x"d4"),
  3137 => (x"49",x"66",x"cc",x"78"),
  3138 => (x"9a",x"ff",x"c3",x"4a"),
  3139 => (x"66",x"cc",x"78",x"72"),
  3140 => (x"c3",x"2a",x"c8",x"4a"),
  3141 => (x"66",x"d0",x"9a",x"ff"),
  3142 => (x"73",x"33",x"c7",x"4b"),
  3143 => (x"71",x"78",x"72",x"b2"),
  3144 => (x"fd",x"49",x"74",x"1e"),
  3145 => (x"ff",x"87",x"dd",x"c5"),
  3146 => (x"78",x"c4",x"48",x"d0"),
  3147 => (x"87",x"f6",x"fc",x"26"),
  3148 => (x"c0",x"1e",x"73",x"1e"),
  3149 => (x"c4",x"4b",x"c0",x"e0"),
  3150 => (x"02",x"bf",x"f2",x"cb"),
  3151 => (x"c4",x"87",x"e7",x"c1"),
  3152 => (x"48",x"bf",x"ef",x"f1"),
  3153 => (x"04",x"a8",x"b7",x"c0"),
  3154 => (x"c4",x"87",x"db",x"c1"),
  3155 => (x"ab",x"bf",x"f6",x"cb"),
  3156 => (x"c4",x"87",x"d3",x"02"),
  3157 => (x"49",x"bf",x"ce",x"cc"),
  3158 => (x"1e",x"71",x"81",x"d0"),
  3159 => (x"49",x"fe",x"cb",x"c4"),
  3160 => (x"87",x"cc",x"e8",x"fd"),
  3161 => (x"1e",x"73",x"86",x"c4"),
  3162 => (x"1e",x"e6",x"cc",x"c4"),
  3163 => (x"49",x"fe",x"cb",x"c4"),
  3164 => (x"87",x"e3",x"e9",x"fd"),
  3165 => (x"cb",x"c4",x"86",x"c8"),
  3166 => (x"02",x"ab",x"bf",x"f6"),
  3167 => (x"c0",x"49",x"87",x"d6"),
  3168 => (x"c4",x"89",x"d0",x"e0"),
  3169 => (x"81",x"bf",x"ce",x"cc"),
  3170 => (x"cb",x"c4",x"1e",x"71"),
  3171 => (x"e7",x"fd",x"49",x"fe"),
  3172 => (x"86",x"c4",x"87",x"de"),
  3173 => (x"1e",x"49",x"66",x"c8"),
  3174 => (x"cc",x"c4",x"1e",x"73"),
  3175 => (x"d1",x"fd",x"49",x"e6"),
  3176 => (x"c0",x"86",x"c8",x"87"),
  3177 => (x"e4",x"c0",x"87",x"e1"),
  3178 => (x"cc",x"c4",x"1e",x"f0"),
  3179 => (x"cb",x"c4",x"1e",x"e6"),
  3180 => (x"e8",x"fd",x"49",x"fe"),
  3181 => (x"66",x"d0",x"87",x"e1"),
  3182 => (x"e4",x"c0",x"1e",x"49"),
  3183 => (x"cc",x"c4",x"1e",x"f0"),
  3184 => (x"ed",x"fc",x"49",x"e6"),
  3185 => (x"fa",x"86",x"d0",x"87"),
  3186 => (x"c4",x"1e",x"87",x"de"),
  3187 => (x"05",x"bf",x"c6",x"cc"),
  3188 => (x"f1",x"c4",x"87",x"db"),
  3189 => (x"50",x"c1",x"48",x"de"),
  3190 => (x"cb",x"1e",x"1e",x"c0"),
  3191 => (x"fb",x"49",x"c2",x"1e"),
  3192 => (x"86",x"cc",x"87",x"c7"),
  3193 => (x"d5",x"fb",x"49",x"c1"),
  3194 => (x"c2",x"48",x"c0",x"87"),
  3195 => (x"26",x"48",x"c1",x"87"),
  3196 => (x"1e",x"73",x"1e",x"4f"),
  3197 => (x"bf",x"da",x"f1",x"c4"),
  3198 => (x"06",x"a8",x"c0",x"48"),
  3199 => (x"c3",x"87",x"e9",x"c0"),
  3200 => (x"49",x"bf",x"d6",x"eb"),
  3201 => (x"87",x"de",x"e3",x"c0"),
  3202 => (x"c7",x"02",x"98",x"70"),
  3203 => (x"49",x"cd",x"87",x"e3"),
  3204 => (x"87",x"c6",x"e3",x"c0"),
  3205 => (x"eb",x"c3",x"49",x"70"),
  3206 => (x"f1",x"c4",x"59",x"da"),
  3207 => (x"c1",x"48",x"bf",x"da"),
  3208 => (x"de",x"f1",x"c4",x"88"),
  3209 => (x"87",x"c9",x"c7",x"58"),
  3210 => (x"97",x"de",x"f1",x"c4"),
  3211 => (x"aa",x"c2",x"4a",x"bf"),
  3212 => (x"87",x"ca",x"c3",x"05"),
  3213 => (x"bf",x"eb",x"f1",x"c4"),
  3214 => (x"de",x"cb",x"c4",x"48"),
  3215 => (x"06",x"a8",x"b7",x"bf"),
  3216 => (x"f1",x"c4",x"87",x"c9"),
  3217 => (x"50",x"c0",x"48",x"de"),
  3218 => (x"c4",x"87",x"e6",x"c6"),
  3219 => (x"bf",x"97",x"e9",x"f1"),
  3220 => (x"87",x"dd",x"c6",x"02"),
  3221 => (x"bf",x"c6",x"cc",x"c4"),
  3222 => (x"c4",x"87",x"da",x"05"),
  3223 => (x"c1",x"48",x"de",x"f1"),
  3224 => (x"1e",x"1e",x"c0",x"50"),
  3225 => (x"49",x"c2",x"1e",x"cb"),
  3226 => (x"cc",x"87",x"fe",x"f8"),
  3227 => (x"f9",x"49",x"c1",x"86"),
  3228 => (x"fc",x"c5",x"87",x"f2"),
  3229 => (x"e9",x"f1",x"c4",x"87"),
  3230 => (x"c4",x"50",x"c0",x"48"),
  3231 => (x"02",x"bf",x"f2",x"cb"),
  3232 => (x"1e",x"c1",x"87",x"cd"),
  3233 => (x"49",x"c0",x"e0",x"c0"),
  3234 => (x"c4",x"87",x"e5",x"fa"),
  3235 => (x"c4",x"87",x"d5",x"86"),
  3236 => (x"48",x"bf",x"ef",x"f1"),
  3237 => (x"bf",x"ea",x"cb",x"c4"),
  3238 => (x"c0",x"04",x"a8",x"b7"),
  3239 => (x"f1",x"c4",x"87",x"c6"),
  3240 => (x"50",x"c0",x"48",x"df"),
  3241 => (x"bf",x"f3",x"f1",x"c4"),
  3242 => (x"c4",x"88",x"c1",x"48"),
  3243 => (x"70",x"58",x"f7",x"f1"),
  3244 => (x"cb",x"c0",x"05",x"98"),
  3245 => (x"f8",x"49",x"c0",x"87"),
  3246 => (x"f1",x"c4",x"87",x"ea"),
  3247 => (x"50",x"c0",x"48",x"de"),
  3248 => (x"bf",x"ef",x"f1",x"c4"),
  3249 => (x"c4",x"80",x"c1",x"48"),
  3250 => (x"c4",x"58",x"f3",x"f1"),
  3251 => (x"b7",x"bf",x"ee",x"cb"),
  3252 => (x"dc",x"c4",x"04",x"a8"),
  3253 => (x"eb",x"f1",x"c4",x"87"),
  3254 => (x"80",x"c1",x"48",x"bf"),
  3255 => (x"58",x"ef",x"f1",x"c4"),
  3256 => (x"e1",x"e1",x"49",x"70"),
  3257 => (x"df",x"f1",x"c4",x"87"),
  3258 => (x"c4",x"50",x"c1",x"48"),
  3259 => (x"49",x"bf",x"e6",x"cb"),
  3260 => (x"fe",x"cb",x"c4",x"1e"),
  3261 => (x"f7",x"e1",x"fd",x"49"),
  3262 => (x"c3",x"86",x"c4",x"87"),
  3263 => (x"aa",x"c3",x"87",x"f3"),
  3264 => (x"87",x"ed",x"c3",x"05"),
  3265 => (x"bf",x"c6",x"cc",x"c4"),
  3266 => (x"87",x"da",x"c0",x"05"),
  3267 => (x"48",x"de",x"f1",x"c4"),
  3268 => (x"1e",x"c0",x"50",x"c1"),
  3269 => (x"c2",x"1e",x"cb",x"1e"),
  3270 => (x"87",x"cd",x"f6",x"49"),
  3271 => (x"49",x"c1",x"86",x"cc"),
  3272 => (x"c3",x"87",x"c1",x"f7"),
  3273 => (x"f1",x"c4",x"87",x"cb"),
  3274 => (x"f2",x"49",x"bf",x"ef"),
  3275 => (x"f1",x"c4",x"87",x"cd"),
  3276 => (x"f1",x"c4",x"58",x"ef"),
  3277 => (x"05",x"bf",x"97",x"ea"),
  3278 => (x"c0",x"87",x"d5",x"c1"),
  3279 => (x"cb",x"f2",x"c4",x"4b"),
  3280 => (x"b7",x"c0",x"48",x"bf"),
  3281 => (x"c7",x"c1",x"04",x"a8"),
  3282 => (x"f2",x"cb",x"c4",x"87"),
  3283 => (x"e8",x"c0",x"05",x"bf"),
  3284 => (x"ef",x"f1",x"c4",x"87"),
  3285 => (x"cb",x"c4",x"49",x"bf"),
  3286 => (x"c0",x"89",x"bf",x"ea"),
  3287 => (x"c4",x"91",x"f0",x"e4"),
  3288 => (x"81",x"bf",x"e6",x"cb"),
  3289 => (x"cb",x"c4",x"1e",x"71"),
  3290 => (x"e0",x"fd",x"49",x"fe"),
  3291 => (x"1e",x"c0",x"87",x"c2"),
  3292 => (x"49",x"f0",x"e4",x"c0"),
  3293 => (x"c8",x"87",x"f9",x"f6"),
  3294 => (x"ef",x"f1",x"c4",x"86"),
  3295 => (x"80",x"c1",x"48",x"bf"),
  3296 => (x"58",x"f3",x"f1",x"c4"),
  3297 => (x"f2",x"c4",x"83",x"c1"),
  3298 => (x"ab",x"b7",x"bf",x"cb"),
  3299 => (x"87",x"f9",x"fe",x"06"),
  3300 => (x"48",x"cb",x"f2",x"c4"),
  3301 => (x"f1",x"c4",x"78",x"c0"),
  3302 => (x"c4",x"48",x"bf",x"ef"),
  3303 => (x"b7",x"bf",x"c7",x"f2"),
  3304 => (x"d7",x"c0",x"03",x"a8"),
  3305 => (x"f2",x"cb",x"c4",x"87"),
  3306 => (x"cf",x"c0",x"05",x"bf"),
  3307 => (x"eb",x"f1",x"c4",x"87"),
  3308 => (x"cb",x"c4",x"48",x"bf"),
  3309 => (x"a8",x"b7",x"bf",x"de"),
  3310 => (x"87",x"f5",x"c0",x"06"),
  3311 => (x"97",x"cf",x"f2",x"c4"),
  3312 => (x"a9",x"c1",x"49",x"bf"),
  3313 => (x"87",x"d2",x"c0",x"05"),
  3314 => (x"48",x"ef",x"f1",x"c4"),
  3315 => (x"bf",x"c3",x"f2",x"c4"),
  3316 => (x"da",x"f1",x"c4",x"78"),
  3317 => (x"c0",x"78",x"c2",x"48"),
  3318 => (x"f1",x"c4",x"87",x"c6"),
  3319 => (x"50",x"c0",x"48",x"de"),
  3320 => (x"97",x"cf",x"f2",x"c4"),
  3321 => (x"a9",x"c2",x"49",x"bf"),
  3322 => (x"87",x"c5",x"c0",x"05"),
  3323 => (x"f3",x"f3",x"49",x"c0"),
  3324 => (x"87",x"f4",x"f1",x"87"),
  3325 => (x"5c",x"5b",x"5e",x"0e"),
  3326 => (x"c4",x"ff",x"0e",x"5d"),
  3327 => (x"c0",x"4b",x"76",x"86"),
  3328 => (x"49",x"e0",x"c0",x"4a"),
  3329 => (x"87",x"ce",x"f3",x"fc"),
  3330 => (x"c8",x"48",x"d0",x"ff"),
  3331 => (x"d4",x"ff",x"78",x"c5"),
  3332 => (x"78",x"e2",x"c1",x"48"),
  3333 => (x"48",x"a6",x"e0",x"c0"),
  3334 => (x"d4",x"ff",x"78",x"c0"),
  3335 => (x"c0",x"78",x"c0",x"48"),
  3336 => (x"c0",x"49",x"a6",x"e4"),
  3337 => (x"68",x"81",x"66",x"e0"),
  3338 => (x"66",x"e0",x"c0",x"51"),
  3339 => (x"c0",x"80",x"c1",x"48"),
  3340 => (x"cc",x"58",x"a6",x"e4"),
  3341 => (x"ff",x"04",x"a8",x"b7"),
  3342 => (x"d0",x"ff",x"87",x"e0"),
  3343 => (x"c0",x"78",x"c4",x"48"),
  3344 => (x"4c",x"66",x"97",x"e4"),
  3345 => (x"f3",x"c0",x"02",x"9c"),
  3346 => (x"02",x"8c",x"c3",x"87"),
  3347 => (x"c5",x"87",x"fe",x"c0"),
  3348 => (x"e5",x"c6",x"02",x"8c"),
  3349 => (x"02",x"8c",x"cd",x"87"),
  3350 => (x"c3",x"87",x"e9",x"c8"),
  3351 => (x"c8",x"02",x"8c",x"c3"),
  3352 => (x"8c",x"c1",x"87",x"fb"),
  3353 => (x"87",x"d2",x"cc",x"02"),
  3354 => (x"c9",x"d0",x"02",x"8c"),
  3355 => (x"02",x"8c",x"c3",x"87"),
  3356 => (x"c1",x"87",x"da",x"d0"),
  3357 => (x"f8",x"c1",x"02",x"8c"),
  3358 => (x"87",x"cc",x"d4",x"87"),
  3359 => (x"70",x"87",x"cb",x"f5"),
  3360 => (x"dd",x"d4",x"02",x"98"),
  3361 => (x"f0",x"49",x"c0",x"87"),
  3362 => (x"d5",x"d4",x"87",x"f4"),
  3363 => (x"7e",x"97",x"d2",x"87"),
  3364 => (x"c2",x"48",x"a6",x"c1"),
  3365 => (x"f0",x"c1",x"50",x"c0"),
  3366 => (x"c4",x"80",x"c1",x"50"),
  3367 => (x"bf",x"97",x"d6",x"f1"),
  3368 => (x"ca",x"80",x"c4",x"50"),
  3369 => (x"c4",x"80",x"c4",x"50"),
  3370 => (x"bf",x"97",x"d7",x"f1"),
  3371 => (x"d8",x"f1",x"c4",x"50"),
  3372 => (x"c4",x"50",x"bf",x"97"),
  3373 => (x"bf",x"97",x"d9",x"f1"),
  3374 => (x"d9",x"f1",x"c4",x"50"),
  3375 => (x"c4",x"50",x"c0",x"48"),
  3376 => (x"c4",x"48",x"d8",x"f1"),
  3377 => (x"bf",x"97",x"d9",x"f1"),
  3378 => (x"d7",x"f1",x"c4",x"50"),
  3379 => (x"d8",x"f1",x"c4",x"48"),
  3380 => (x"c4",x"50",x"bf",x"97"),
  3381 => (x"c4",x"48",x"d6",x"f1"),
  3382 => (x"bf",x"97",x"d7",x"f1"),
  3383 => (x"d2",x"1e",x"c1",x"50"),
  3384 => (x"49",x"a6",x"ca",x"1e"),
  3385 => (x"c8",x"87",x"cb",x"f0"),
  3386 => (x"ef",x"49",x"c0",x"86"),
  3387 => (x"f1",x"d2",x"87",x"d0"),
  3388 => (x"87",x"d6",x"f3",x"87"),
  3389 => (x"d2",x"02",x"98",x"70"),
  3390 => (x"e5",x"c0",x"87",x"e8"),
  3391 => (x"c0",x"48",x"66",x"97"),
  3392 => (x"70",x"58",x"a6",x"e4"),
  3393 => (x"87",x"da",x"02",x"98"),
  3394 => (x"c0",x"88",x"c1",x"48"),
  3395 => (x"70",x"58",x"a6",x"e4"),
  3396 => (x"ed",x"c0",x"02",x"98"),
  3397 => (x"88",x"c1",x"48",x"87"),
  3398 => (x"58",x"a6",x"e4",x"c0"),
  3399 => (x"c1",x"02",x"98",x"70"),
  3400 => (x"97",x"c2",x"87",x"eb"),
  3401 => (x"48",x"a6",x"c1",x"7e"),
  3402 => (x"c1",x"50",x"c0",x"c2"),
  3403 => (x"de",x"cb",x"c4",x"50"),
  3404 => (x"c2",x"ec",x"49",x"bf"),
  3405 => (x"08",x"a6",x"c3",x"87"),
  3406 => (x"a6",x"e0",x"c0",x"50"),
  3407 => (x"c2",x"78",x"c2",x"48"),
  3408 => (x"cb",x"c4",x"87",x"e2"),
  3409 => (x"c2",x"49",x"bf",x"da"),
  3410 => (x"f0",x"c0",x"81",x"d6"),
  3411 => (x"ff",x"71",x"1e",x"a6"),
  3412 => (x"c4",x"87",x"fd",x"ca"),
  3413 => (x"c1",x"7e",x"97",x"86"),
  3414 => (x"c0",x"c2",x"48",x"a6"),
  3415 => (x"97",x"f0",x"c0",x"50"),
  3416 => (x"d2",x"eb",x"49",x"66"),
  3417 => (x"08",x"a6",x"c2",x"87"),
  3418 => (x"97",x"f1",x"c0",x"50"),
  3419 => (x"c6",x"eb",x"49",x"66"),
  3420 => (x"08",x"a6",x"c3",x"87"),
  3421 => (x"97",x"f2",x"c0",x"50"),
  3422 => (x"fa",x"ea",x"49",x"66"),
  3423 => (x"08",x"a6",x"c4",x"87"),
  3424 => (x"48",x"a6",x"c5",x"50"),
  3425 => (x"80",x"da",x"50",x"c0"),
  3426 => (x"d7",x"c1",x"78",x"c4"),
  3427 => (x"97",x"e6",x"c0",x"87"),
  3428 => (x"ef",x"eb",x"49",x"66"),
  3429 => (x"ea",x"cb",x"c4",x"87"),
  3430 => (x"d6",x"c2",x"49",x"bf"),
  3431 => (x"a6",x"f0",x"c0",x"81"),
  3432 => (x"c9",x"ff",x"71",x"1e"),
  3433 => (x"86",x"c4",x"87",x"ea"),
  3434 => (x"a6",x"c1",x"7e",x"97"),
  3435 => (x"50",x"c0",x"c2",x"48"),
  3436 => (x"66",x"97",x"f0",x"c0"),
  3437 => (x"87",x"ff",x"e9",x"49"),
  3438 => (x"50",x"08",x"a6",x"c2"),
  3439 => (x"66",x"97",x"f1",x"c0"),
  3440 => (x"87",x"f3",x"e9",x"49"),
  3441 => (x"50",x"08",x"a6",x"c3"),
  3442 => (x"66",x"97",x"f2",x"c0"),
  3443 => (x"87",x"e7",x"e9",x"49"),
  3444 => (x"50",x"08",x"a6",x"c4"),
  3445 => (x"bf",x"f2",x"cb",x"c4"),
  3446 => (x"c9",x"31",x"c2",x"49"),
  3447 => (x"48",x"59",x"97",x"a6"),
  3448 => (x"78",x"c4",x"80",x"db"),
  3449 => (x"e4",x"c0",x"1e",x"c1"),
  3450 => (x"a6",x"ca",x"1e",x"66"),
  3451 => (x"87",x"c2",x"ec",x"49"),
  3452 => (x"49",x"c0",x"86",x"c8"),
  3453 => (x"ce",x"87",x"c7",x"eb"),
  3454 => (x"cd",x"ef",x"87",x"e8"),
  3455 => (x"02",x"98",x"70",x"87"),
  3456 => (x"c0",x"87",x"df",x"ce"),
  3457 => (x"49",x"66",x"97",x"e5"),
  3458 => (x"e6",x"c0",x"31",x"d0"),
  3459 => (x"c8",x"4a",x"66",x"97"),
  3460 => (x"c0",x"b1",x"72",x"32"),
  3461 => (x"4a",x"66",x"97",x"e7"),
  3462 => (x"c7",x"4d",x"71",x"b1"),
  3463 => (x"9d",x"ff",x"ff",x"ff"),
  3464 => (x"66",x"97",x"e8",x"c0"),
  3465 => (x"87",x"c8",x"c0",x"02"),
  3466 => (x"a6",x"e4",x"c0",x"48"),
  3467 => (x"87",x"c7",x"c0",x"58"),
  3468 => (x"48",x"a6",x"e0",x"c0"),
  3469 => (x"75",x"78",x"c0",x"c4"),
  3470 => (x"87",x"ff",x"e5",x"49"),
  3471 => (x"58",x"ef",x"f1",x"c4"),
  3472 => (x"48",x"da",x"f1",x"c4"),
  3473 => (x"f1",x"c4",x"78",x"c0"),
  3474 => (x"f1",x"c4",x"5d",x"f3"),
  3475 => (x"e0",x"c0",x"48",x"f3"),
  3476 => (x"49",x"75",x"78",x"66"),
  3477 => (x"bf",x"ea",x"cb",x"c4"),
  3478 => (x"f6",x"cb",x"c4",x"89"),
  3479 => (x"cb",x"c4",x"91",x"bf"),
  3480 => (x"71",x"81",x"bf",x"e6"),
  3481 => (x"fe",x"cb",x"c4",x"1e"),
  3482 => (x"c3",x"d4",x"fd",x"49"),
  3483 => (x"c4",x"86",x"c4",x"87"),
  3484 => (x"c0",x"48",x"ff",x"f1"),
  3485 => (x"e9",x"f1",x"c4",x"78"),
  3486 => (x"c4",x"50",x"c1",x"48"),
  3487 => (x"c2",x"48",x"de",x"f1"),
  3488 => (x"87",x"de",x"cc",x"50"),
  3489 => (x"66",x"97",x"e8",x"c0"),
  3490 => (x"87",x"c9",x"c0",x"02"),
  3491 => (x"48",x"e8",x"f1",x"c4"),
  3492 => (x"cd",x"cc",x"50",x"c1"),
  3493 => (x"e8",x"49",x"c0",x"87"),
  3494 => (x"c5",x"cc",x"87",x"e4"),
  3495 => (x"87",x"ea",x"ec",x"87"),
  3496 => (x"cb",x"02",x"98",x"70"),
  3497 => (x"ed",x"c0",x"87",x"fc"),
  3498 => (x"48",x"49",x"66",x"97"),
  3499 => (x"c0",x"98",x"c0",x"c3"),
  3500 => (x"70",x"58",x"a6",x"e4"),
  3501 => (x"dc",x"c0",x"02",x"98"),
  3502 => (x"c0",x"c1",x"48",x"87"),
  3503 => (x"a6",x"e4",x"c0",x"88"),
  3504 => (x"02",x"98",x"70",x"58"),
  3505 => (x"48",x"87",x"e9",x"c0"),
  3506 => (x"c0",x"88",x"c0",x"c1"),
  3507 => (x"70",x"58",x"a6",x"e4"),
  3508 => (x"c7",x"c1",x"02",x"98"),
  3509 => (x"97",x"e7",x"c0",x"87"),
  3510 => (x"31",x"d0",x"49",x"66"),
  3511 => (x"66",x"97",x"e8",x"c0"),
  3512 => (x"72",x"32",x"c8",x"4a"),
  3513 => (x"97",x"e9",x"c0",x"b1"),
  3514 => (x"71",x"4d",x"4a",x"66"),
  3515 => (x"87",x"f9",x"c0",x"b5"),
  3516 => (x"66",x"97",x"e8",x"c0"),
  3517 => (x"87",x"f4",x"e5",x"49"),
  3518 => (x"c0",x"1e",x"49",x"70"),
  3519 => (x"49",x"66",x"97",x"eb"),
  3520 => (x"70",x"87",x"e9",x"e5"),
  3521 => (x"ee",x"c0",x"1e",x"49"),
  3522 => (x"e5",x"49",x"66",x"97"),
  3523 => (x"4a",x"70",x"87",x"de"),
  3524 => (x"cb",x"c5",x"ff",x"49"),
  3525 => (x"70",x"86",x"c8",x"87"),
  3526 => (x"87",x"cd",x"c0",x"4d"),
  3527 => (x"66",x"97",x"e6",x"c0"),
  3528 => (x"87",x"e0",x"e5",x"49"),
  3529 => (x"bf",x"ea",x"cb",x"c4"),
  3530 => (x"da",x"f1",x"c4",x"4d"),
  3531 => (x"c4",x"78",x"c0",x"48"),
  3532 => (x"75",x"5d",x"f3",x"f1"),
  3533 => (x"87",x"c3",x"e2",x"49"),
  3534 => (x"58",x"ef",x"f1",x"c4"),
  3535 => (x"5d",x"c7",x"f2",x"c4"),
  3536 => (x"48",x"c7",x"f2",x"c4"),
  3537 => (x"bf",x"da",x"cb",x"c4"),
  3538 => (x"cf",x"f2",x"c4",x"78"),
  3539 => (x"97",x"e5",x"c0",x"48"),
  3540 => (x"f2",x"c4",x"50",x"66"),
  3541 => (x"78",x"c1",x"48",x"cb"),
  3542 => (x"97",x"cf",x"f2",x"c4"),
  3543 => (x"05",x"99",x"49",x"bf"),
  3544 => (x"c4",x"87",x"c9",x"c0"),
  3545 => (x"c4",x"48",x"de",x"f1"),
  3546 => (x"87",x"c6",x"c0",x"50"),
  3547 => (x"48",x"de",x"f1",x"c4"),
  3548 => (x"49",x"c0",x"50",x"c3"),
  3549 => (x"c8",x"87",x"ed",x"e5"),
  3550 => (x"cd",x"e9",x"87",x"e8"),
  3551 => (x"02",x"98",x"70",x"87"),
  3552 => (x"c0",x"87",x"df",x"c8"),
  3553 => (x"49",x"66",x"97",x"ed"),
  3554 => (x"98",x"c0",x"c3",x"48"),
  3555 => (x"58",x"a6",x"e4",x"c0"),
  3556 => (x"c0",x"02",x"98",x"70"),
  3557 => (x"c1",x"48",x"87",x"dc"),
  3558 => (x"e4",x"c0",x"88",x"c0"),
  3559 => (x"98",x"70",x"58",x"a6"),
  3560 => (x"87",x"e9",x"c0",x"02"),
  3561 => (x"88",x"c0",x"c1",x"48"),
  3562 => (x"58",x"a6",x"e4",x"c0"),
  3563 => (x"c1",x"02",x"98",x"70"),
  3564 => (x"e7",x"c0",x"87",x"c7"),
  3565 => (x"d0",x"49",x"66",x"97"),
  3566 => (x"97",x"e8",x"c0",x"31"),
  3567 => (x"32",x"c8",x"4a",x"66"),
  3568 => (x"e9",x"c0",x"b1",x"72"),
  3569 => (x"4d",x"4a",x"66",x"97"),
  3570 => (x"ee",x"c1",x"b5",x"71"),
  3571 => (x"97",x"e8",x"c0",x"87"),
  3572 => (x"d7",x"e2",x"49",x"66"),
  3573 => (x"1e",x"49",x"70",x"87"),
  3574 => (x"66",x"97",x"eb",x"c0"),
  3575 => (x"87",x"cc",x"e2",x"49"),
  3576 => (x"c0",x"1e",x"49",x"70"),
  3577 => (x"49",x"66",x"97",x"ee"),
  3578 => (x"70",x"87",x"c1",x"e2"),
  3579 => (x"c1",x"ff",x"49",x"4a"),
  3580 => (x"86",x"c8",x"87",x"ee"),
  3581 => (x"c2",x"c1",x"4d",x"70"),
  3582 => (x"97",x"e6",x"c0",x"87"),
  3583 => (x"eb",x"e1",x"49",x"66"),
  3584 => (x"48",x"49",x"70",x"87"),
  3585 => (x"58",x"a6",x"e4",x"c0"),
  3586 => (x"c0",x"05",x"98",x"70"),
  3587 => (x"e0",x"c0",x"87",x"c6"),
  3588 => (x"78",x"c1",x"48",x"a6"),
  3589 => (x"48",x"66",x"e0",x"c0"),
  3590 => (x"bf",x"de",x"cb",x"c4"),
  3591 => (x"c0",x"06",x"a8",x"b7"),
  3592 => (x"e0",x"c0",x"87",x"cc"),
  3593 => (x"cb",x"c4",x"48",x"a6"),
  3594 => (x"c0",x"78",x"bf",x"da"),
  3595 => (x"e0",x"c0",x"87",x"c9"),
  3596 => (x"cb",x"c4",x"48",x"a6"),
  3597 => (x"c0",x"78",x"bf",x"ee"),
  3598 => (x"c4",x"4d",x"66",x"e0"),
  3599 => (x"c0",x"48",x"cf",x"f2"),
  3600 => (x"50",x"66",x"97",x"e5"),
  3601 => (x"5d",x"cb",x"f2",x"c4"),
  3602 => (x"97",x"cf",x"f2",x"c4"),
  3603 => (x"05",x"99",x"49",x"bf"),
  3604 => (x"c4",x"87",x"c9",x"c0"),
  3605 => (x"c0",x"48",x"de",x"f1"),
  3606 => (x"87",x"c6",x"c0",x"50"),
  3607 => (x"48",x"de",x"f1",x"c4"),
  3608 => (x"f2",x"c4",x"50",x"c3"),
  3609 => (x"49",x"bf",x"97",x"cf"),
  3610 => (x"c4",x"02",x"a9",x"c2"),
  3611 => (x"49",x"c0",x"87",x"f4"),
  3612 => (x"c4",x"87",x"cb",x"e1"),
  3613 => (x"d1",x"e5",x"87",x"ec"),
  3614 => (x"02",x"98",x"70",x"87"),
  3615 => (x"c4",x"87",x"e3",x"c4"),
  3616 => (x"c4",x"48",x"de",x"f1"),
  3617 => (x"e0",x"49",x"c0",x"50"),
  3618 => (x"d5",x"c4",x"87",x"f4"),
  3619 => (x"87",x"fa",x"e4",x"87"),
  3620 => (x"c4",x"02",x"98",x"70"),
  3621 => (x"f1",x"c4",x"87",x"cc"),
  3622 => (x"c4",x"48",x"bf",x"ef"),
  3623 => (x"88",x"bf",x"ea",x"cb"),
  3624 => (x"58",x"a6",x"e4",x"c0"),
  3625 => (x"c1",x"7e",x"97",x"ca"),
  3626 => (x"c0",x"c2",x"48",x"a6"),
  3627 => (x"de",x"f1",x"c4",x"50"),
  3628 => (x"c0",x"48",x"bf",x"97"),
  3629 => (x"c4",x"58",x"a6",x"f7"),
  3630 => (x"c9",x"c0",x"05",x"a8"),
  3631 => (x"a6",x"f3",x"c0",x"87"),
  3632 => (x"c0",x"78",x"c2",x"48"),
  3633 => (x"f3",x"c0",x"87",x"e1"),
  3634 => (x"a8",x"c3",x"48",x"66"),
  3635 => (x"87",x"c9",x"c0",x"05"),
  3636 => (x"48",x"a6",x"f7",x"c0"),
  3637 => (x"c6",x"c0",x"78",x"c0"),
  3638 => (x"a6",x"f7",x"c0",x"87"),
  3639 => (x"c0",x"78",x"c3",x"48"),
  3640 => (x"c0",x"48",x"a6",x"f3"),
  3641 => (x"c2",x"78",x"66",x"f7"),
  3642 => (x"f3",x"c0",x"48",x"a6"),
  3643 => (x"50",x"c0",x"50",x"66"),
  3644 => (x"bf",x"eb",x"f1",x"c4"),
  3645 => (x"ff",x"81",x"c1",x"49"),
  3646 => (x"c4",x"87",x"fc",x"dc"),
  3647 => (x"c4",x"50",x"08",x"a6"),
  3648 => (x"49",x"bf",x"eb",x"f1"),
  3649 => (x"87",x"ef",x"dc",x"ff"),
  3650 => (x"50",x"08",x"a6",x"c5"),
  3651 => (x"4b",x"a6",x"f0",x"c0"),
  3652 => (x"66",x"e4",x"c0",x"1e"),
  3653 => (x"f7",x"fb",x"fe",x"49"),
  3654 => (x"97",x"f4",x"c0",x"87"),
  3655 => (x"dc",x"ff",x"49",x"66"),
  3656 => (x"a6",x"ca",x"87",x"d5"),
  3657 => (x"f5",x"c0",x"50",x"08"),
  3658 => (x"ff",x"49",x"66",x"97"),
  3659 => (x"cb",x"87",x"c8",x"dc"),
  3660 => (x"c0",x"50",x"08",x"a6"),
  3661 => (x"49",x"66",x"97",x"f6"),
  3662 => (x"87",x"fb",x"db",x"ff"),
  3663 => (x"50",x"08",x"a6",x"cc"),
  3664 => (x"f1",x"c4",x"1e",x"73"),
  3665 => (x"fe",x"49",x"bf",x"ef"),
  3666 => (x"c0",x"87",x"c5",x"fb"),
  3667 => (x"49",x"66",x"97",x"f8"),
  3668 => (x"87",x"e3",x"db",x"ff"),
  3669 => (x"50",x"08",x"a6",x"d1"),
  3670 => (x"66",x"97",x"f9",x"c0"),
  3671 => (x"d6",x"db",x"ff",x"49"),
  3672 => (x"08",x"a6",x"d2",x"87"),
  3673 => (x"97",x"fa",x"c0",x"50"),
  3674 => (x"db",x"ff",x"49",x"66"),
  3675 => (x"a6",x"d3",x"87",x"c9"),
  3676 => (x"1e",x"c1",x"50",x"08"),
  3677 => (x"a6",x"d2",x"1e",x"ca"),
  3678 => (x"f5",x"dd",x"ff",x"49"),
  3679 => (x"c0",x"86",x"d0",x"87"),
  3680 => (x"f9",x"dc",x"ff",x"49"),
  3681 => (x"87",x"da",x"c0",x"87"),
  3682 => (x"c0",x"1e",x"1e",x"c0"),
  3683 => (x"49",x"c5",x"1e",x"e0"),
  3684 => (x"87",x"d5",x"dc",x"ff"),
  3685 => (x"f1",x"c4",x"86",x"cc"),
  3686 => (x"78",x"c0",x"48",x"e4"),
  3687 => (x"dc",x"ff",x"49",x"c1"),
  3688 => (x"c4",x"ff",x"87",x"dc"),
  3689 => (x"fb",x"da",x"ff",x"8e"),
  3690 => (x"86",x"f4",x"1e",x"87"),
  3691 => (x"c8",x"48",x"d0",x"ff"),
  3692 => (x"d4",x"ff",x"78",x"c5"),
  3693 => (x"78",x"e3",x"c1",x"48"),
  3694 => (x"d4",x"ff",x"4a",x"c0"),
  3695 => (x"76",x"78",x"c0",x"48"),
  3696 => (x"68",x"81",x"72",x"49"),
  3697 => (x"ca",x"82",x"c1",x"51"),
  3698 => (x"ed",x"04",x"aa",x"b7"),
  3699 => (x"48",x"d0",x"ff",x"87"),
  3700 => (x"8e",x"f4",x"78",x"c4"),
  3701 => (x"c4",x"1e",x"4f",x"26"),
  3702 => (x"c1",x"48",x"e9",x"f1"),
  3703 => (x"1e",x"4f",x"26",x"50"),
  3704 => (x"48",x"da",x"f1",x"c4"),
  3705 => (x"f1",x"c4",x"78",x"c0"),
  3706 => (x"40",x"c0",x"48",x"eb"),
  3707 => (x"f7",x"f1",x"c4",x"78"),
  3708 => (x"c4",x"78",x"c0",x"48"),
  3709 => (x"c1",x"48",x"df",x"f1"),
  3710 => (x"c6",x"cc",x"c4",x"50"),
  3711 => (x"87",x"c4",x"02",x"bf"),
  3712 => (x"87",x"c2",x"49",x"c0"),
  3713 => (x"f1",x"c4",x"49",x"c1"),
  3714 => (x"c4",x"59",x"97",x"e2"),
  3715 => (x"c0",x"48",x"fb",x"f1"),
  3716 => (x"f1",x"c4",x"78",x"40"),
  3717 => (x"40",x"c0",x"48",x"e4"),
  3718 => (x"f2",x"c4",x"50",x"50"),
  3719 => (x"40",x"c0",x"48",x"c3"),
  3720 => (x"cf",x"f2",x"c4",x"78"),
  3721 => (x"9f",x"50",x"c0",x"48"),
  3722 => (x"ea",x"f1",x"c4",x"78"),
  3723 => (x"26",x"50",x"c1",x"48"),
  3724 => (x"1e",x"73",x"1e",x"4f"),
  3725 => (x"c8",x"48",x"d0",x"ff"),
  3726 => (x"d4",x"ff",x"78",x"c5"),
  3727 => (x"78",x"e0",x"c1",x"48"),
  3728 => (x"ff",x"c3",x"49",x"68"),
  3729 => (x"48",x"d0",x"ff",x"99"),
  3730 => (x"4b",x"71",x"78",x"c4"),
  3731 => (x"02",x"99",x"c1",x"49"),
  3732 => (x"df",x"e6",x"87",x"c3"),
  3733 => (x"c2",x"49",x"73",x"87"),
  3734 => (x"87",x"c3",x"02",x"99"),
  3735 => (x"73",x"87",x"ca",x"fd"),
  3736 => (x"02",x"99",x"c4",x"49"),
  3737 => (x"ed",x"fd",x"87",x"c3"),
  3738 => (x"c8",x"49",x"73",x"87"),
  3739 => (x"87",x"d6",x"02",x"99"),
  3740 => (x"ff",x"87",x"ec",x"fd"),
  3741 => (x"c5",x"c8",x"48",x"d0"),
  3742 => (x"48",x"d4",x"ff",x"78"),
  3743 => (x"c0",x"78",x"e6",x"c1"),
  3744 => (x"48",x"d0",x"ff",x"78"),
  3745 => (x"49",x"73",x"78",x"c4"),
  3746 => (x"f1",x"c4",x"99",x"d0"),
  3747 => (x"ff",x"59",x"97",x"ee"),
  3748 => (x"c4",x"87",x"de",x"dd"),
  3749 => (x"02",x"bf",x"e4",x"f1"),
  3750 => (x"f1",x"c4",x"87",x"d7"),
  3751 => (x"d0",x"05",x"bf",x"da"),
  3752 => (x"d0",x"f2",x"c4",x"87"),
  3753 => (x"ff",x"49",x"bf",x"9f"),
  3754 => (x"c4",x"87",x"d3",x"d8"),
  3755 => (x"c0",x"48",x"e4",x"f1"),
  3756 => (x"e8",x"f1",x"c4",x"78"),
  3757 => (x"d9",x"02",x"bf",x"97"),
  3758 => (x"48",x"d0",x"ff",x"87"),
  3759 => (x"ff",x"78",x"c5",x"c8"),
  3760 => (x"e5",x"c1",x"48",x"d4"),
  3761 => (x"ff",x"78",x"c0",x"78"),
  3762 => (x"78",x"c4",x"48",x"d0"),
  3763 => (x"48",x"e8",x"f1",x"c4"),
  3764 => (x"d6",x"ff",x"50",x"c0"),
  3765 => (x"00",x"00",x"87",x"d2"),
  3766 => (x"71",x"1e",x"00",x"00"),
  3767 => (x"bf",x"c8",x"ff",x"4a"),
  3768 => (x"48",x"a1",x"72",x"49"),
  3769 => (x"ff",x"1e",x"4f",x"26"),
  3770 => (x"fe",x"89",x"bf",x"c8"),
  3771 => (x"c0",x"c0",x"c0",x"c0"),
  3772 => (x"c4",x"01",x"a9",x"c0"),
  3773 => (x"c2",x"4a",x"c0",x"87"),
  3774 => (x"72",x"4a",x"c1",x"87"),
  3775 => (x"0e",x"4f",x"26",x"48"),
  3776 => (x"5d",x"5c",x"5b",x"5e"),
  3777 => (x"ff",x"4b",x"71",x"0e"),
  3778 => (x"66",x"d0",x"4c",x"d4"),
  3779 => (x"d6",x"78",x"c0",x"48"),
  3780 => (x"df",x"cf",x"fe",x"49"),
  3781 => (x"7c",x"ff",x"c3",x"87"),
  3782 => (x"ff",x"c3",x"49",x"6c"),
  3783 => (x"49",x"4d",x"71",x"99"),
  3784 => (x"c1",x"99",x"f0",x"c3"),
  3785 => (x"cb",x"05",x"a9",x"e0"),
  3786 => (x"7c",x"ff",x"c3",x"87"),
  3787 => (x"98",x"c3",x"48",x"6c"),
  3788 => (x"78",x"08",x"66",x"d0"),
  3789 => (x"6c",x"7c",x"ff",x"c3"),
  3790 => (x"31",x"c8",x"49",x"4a"),
  3791 => (x"6c",x"7c",x"ff",x"c3"),
  3792 => (x"72",x"b2",x"71",x"4a"),
  3793 => (x"c3",x"31",x"c8",x"49"),
  3794 => (x"4a",x"6c",x"7c",x"ff"),
  3795 => (x"49",x"72",x"b2",x"71"),
  3796 => (x"ff",x"c3",x"31",x"c8"),
  3797 => (x"71",x"4a",x"6c",x"7c"),
  3798 => (x"48",x"d0",x"ff",x"b2"),
  3799 => (x"73",x"78",x"e0",x"c0"),
  3800 => (x"87",x"c2",x"02",x"9b"),
  3801 => (x"48",x"75",x"7b",x"72"),
  3802 => (x"4c",x"26",x"4d",x"26"),
  3803 => (x"4f",x"26",x"4b",x"26"),
  3804 => (x"0e",x"4f",x"26",x"1e"),
  3805 => (x"0e",x"5c",x"5b",x"5e"),
  3806 => (x"1e",x"76",x"86",x"f8"),
  3807 => (x"fd",x"49",x"a6",x"c8"),
  3808 => (x"86",x"c4",x"87",x"fd"),
  3809 => (x"48",x"6e",x"4b",x"70"),
  3810 => (x"c2",x"01",x"a8",x"c0"),
  3811 => (x"4a",x"73",x"87",x"f0"),
  3812 => (x"c1",x"9a",x"f0",x"c3"),
  3813 => (x"c7",x"02",x"aa",x"d0"),
  3814 => (x"aa",x"e0",x"c1",x"87"),
  3815 => (x"87",x"de",x"c2",x"05"),
  3816 => (x"99",x"c8",x"49",x"73"),
  3817 => (x"ff",x"87",x"c3",x"02"),
  3818 => (x"4c",x"73",x"87",x"c6"),
  3819 => (x"ac",x"c2",x"9c",x"c3"),
  3820 => (x"87",x"c2",x"c1",x"05"),
  3821 => (x"c9",x"49",x"66",x"c4"),
  3822 => (x"c4",x"1e",x"71",x"31"),
  3823 => (x"92",x"d4",x"4a",x"66"),
  3824 => (x"49",x"d2",x"f2",x"c4"),
  3825 => (x"fe",x"fc",x"81",x"72"),
  3826 => (x"49",x"d8",x"87",x"e6"),
  3827 => (x"87",x"e4",x"cc",x"fe"),
  3828 => (x"c3",x"1e",x"c0",x"c8"),
  3829 => (x"fc",x"49",x"ca",x"fa"),
  3830 => (x"ff",x"87",x"ff",x"da"),
  3831 => (x"e0",x"c0",x"48",x"d0"),
  3832 => (x"ca",x"fa",x"c3",x"78"),
  3833 => (x"4a",x"66",x"cc",x"1e"),
  3834 => (x"f2",x"c4",x"92",x"d4"),
  3835 => (x"81",x"72",x"49",x"d2"),
  3836 => (x"87",x"f9",x"fc",x"fc"),
  3837 => (x"ac",x"c1",x"86",x"cc"),
  3838 => (x"87",x"c2",x"c1",x"05"),
  3839 => (x"c9",x"49",x"66",x"c4"),
  3840 => (x"c4",x"1e",x"71",x"31"),
  3841 => (x"92",x"d4",x"4a",x"66"),
  3842 => (x"49",x"d2",x"f2",x"c4"),
  3843 => (x"fd",x"fc",x"81",x"72"),
  3844 => (x"fa",x"c3",x"87",x"de"),
  3845 => (x"66",x"c8",x"1e",x"ca"),
  3846 => (x"c4",x"92",x"d4",x"4a"),
  3847 => (x"72",x"49",x"d2",x"f2"),
  3848 => (x"c5",x"fb",x"fc",x"81"),
  3849 => (x"fe",x"49",x"d7",x"87"),
  3850 => (x"c8",x"87",x"c9",x"cb"),
  3851 => (x"fa",x"c3",x"1e",x"c0"),
  3852 => (x"d9",x"fc",x"49",x"ca"),
  3853 => (x"86",x"cc",x"87",x"ce"),
  3854 => (x"c0",x"48",x"d0",x"ff"),
  3855 => (x"8e",x"f8",x"78",x"e0"),
  3856 => (x"0e",x"87",x"e7",x"fc"),
  3857 => (x"5d",x"5c",x"5b",x"5e"),
  3858 => (x"4d",x"71",x"1e",x"0e"),
  3859 => (x"d4",x"4c",x"d4",x"ff"),
  3860 => (x"c3",x"48",x"7e",x"66"),
  3861 => (x"c5",x"06",x"a8",x"b7"),
  3862 => (x"c1",x"48",x"c0",x"87"),
  3863 => (x"49",x"75",x"87",x"e2"),
  3864 => (x"87",x"ca",x"d1",x"fd"),
  3865 => (x"66",x"c4",x"1e",x"75"),
  3866 => (x"c4",x"93",x"d4",x"4b"),
  3867 => (x"73",x"83",x"d2",x"f2"),
  3868 => (x"d9",x"f6",x"fc",x"49"),
  3869 => (x"6b",x"83",x"c8",x"87"),
  3870 => (x"48",x"d0",x"ff",x"4b"),
  3871 => (x"dd",x"78",x"e1",x"c8"),
  3872 => (x"c3",x"49",x"73",x"7c"),
  3873 => (x"7c",x"71",x"99",x"ff"),
  3874 => (x"b7",x"c8",x"49",x"73"),
  3875 => (x"99",x"ff",x"c3",x"29"),
  3876 => (x"49",x"73",x"7c",x"71"),
  3877 => (x"c3",x"29",x"b7",x"d0"),
  3878 => (x"7c",x"71",x"99",x"ff"),
  3879 => (x"b7",x"d8",x"49",x"73"),
  3880 => (x"c0",x"7c",x"71",x"29"),
  3881 => (x"7c",x"7c",x"7c",x"7c"),
  3882 => (x"7c",x"7c",x"7c",x"7c"),
  3883 => (x"7c",x"7c",x"7c",x"7c"),
  3884 => (x"c4",x"78",x"e0",x"c0"),
  3885 => (x"49",x"dc",x"1e",x"66"),
  3886 => (x"87",x"dd",x"c9",x"fe"),
  3887 => (x"48",x"73",x"86",x"c8"),
  3888 => (x"87",x"e4",x"fa",x"26"),
  3889 => (x"5c",x"5b",x"5e",x"0e"),
  3890 => (x"71",x"1e",x"0e",x"5d"),
  3891 => (x"4b",x"d4",x"ff",x"7e"),
  3892 => (x"f2",x"c4",x"1e",x"6e"),
  3893 => (x"f4",x"fc",x"49",x"e6"),
  3894 => (x"86",x"c4",x"87",x"f4"),
  3895 => (x"02",x"9d",x"4d",x"70"),
  3896 => (x"c4",x"87",x"c3",x"c3"),
  3897 => (x"4c",x"bf",x"ee",x"f2"),
  3898 => (x"cf",x"fd",x"49",x"6e"),
  3899 => (x"d0",x"ff",x"87",x"c0"),
  3900 => (x"78",x"c5",x"c8",x"48"),
  3901 => (x"c0",x"7b",x"d6",x"c1"),
  3902 => (x"c1",x"7b",x"15",x"4a"),
  3903 => (x"b7",x"e0",x"c0",x"82"),
  3904 => (x"87",x"f5",x"04",x"aa"),
  3905 => (x"c4",x"48",x"d0",x"ff"),
  3906 => (x"78",x"c5",x"c8",x"78"),
  3907 => (x"c1",x"7b",x"d3",x"c1"),
  3908 => (x"74",x"78",x"c4",x"7b"),
  3909 => (x"fc",x"c1",x"02",x"9c"),
  3910 => (x"ca",x"fa",x"c3",x"87"),
  3911 => (x"4d",x"c0",x"c8",x"7e"),
  3912 => (x"ac",x"b7",x"c0",x"8c"),
  3913 => (x"c8",x"87",x"c6",x"03"),
  3914 => (x"c0",x"4d",x"a4",x"c0"),
  3915 => (x"fb",x"c6",x"c4",x"4c"),
  3916 => (x"d0",x"49",x"bf",x"97"),
  3917 => (x"87",x"d2",x"02",x"99"),
  3918 => (x"f2",x"c4",x"1e",x"c0"),
  3919 => (x"f6",x"fc",x"49",x"e6"),
  3920 => (x"86",x"c4",x"87",x"e8"),
  3921 => (x"c0",x"4a",x"49",x"70"),
  3922 => (x"fa",x"c3",x"87",x"ef"),
  3923 => (x"f2",x"c4",x"1e",x"ca"),
  3924 => (x"f6",x"fc",x"49",x"e6"),
  3925 => (x"86",x"c4",x"87",x"d4"),
  3926 => (x"ff",x"4a",x"49",x"70"),
  3927 => (x"c5",x"c8",x"48",x"d0"),
  3928 => (x"7b",x"d4",x"c1",x"78"),
  3929 => (x"7b",x"bf",x"97",x"6e"),
  3930 => (x"80",x"c1",x"48",x"6e"),
  3931 => (x"8d",x"c1",x"7e",x"70"),
  3932 => (x"87",x"f0",x"ff",x"05"),
  3933 => (x"c4",x"48",x"d0",x"ff"),
  3934 => (x"05",x"9a",x"72",x"78"),
  3935 => (x"48",x"c0",x"87",x"c5"),
  3936 => (x"c1",x"87",x"e5",x"c0"),
  3937 => (x"e6",x"f2",x"c4",x"1e"),
  3938 => (x"fc",x"f3",x"fc",x"49"),
  3939 => (x"74",x"86",x"c4",x"87"),
  3940 => (x"c4",x"fe",x"05",x"9c"),
  3941 => (x"48",x"d0",x"ff",x"87"),
  3942 => (x"c1",x"78",x"c5",x"c8"),
  3943 => (x"7b",x"c0",x"7b",x"d3"),
  3944 => (x"48",x"c1",x"78",x"c4"),
  3945 => (x"48",x"c0",x"87",x"c2"),
  3946 => (x"26",x"4d",x"26",x"26"),
  3947 => (x"26",x"4b",x"26",x"4c"),
  3948 => (x"5b",x"5e",x"0e",x"4f"),
  3949 => (x"4b",x"71",x"0e",x"5c"),
  3950 => (x"dd",x"02",x"66",x"cc"),
  3951 => (x"f0",x"c0",x"4c",x"87"),
  3952 => (x"87",x"dd",x"02",x"8c"),
  3953 => (x"8a",x"c1",x"4a",x"74"),
  3954 => (x"8a",x"87",x"d6",x"02"),
  3955 => (x"8a",x"87",x"d2",x"02"),
  3956 => (x"d0",x"87",x"ce",x"02"),
  3957 => (x"87",x"db",x"02",x"8a"),
  3958 => (x"49",x"73",x"87",x"df"),
  3959 => (x"d8",x"87",x"e5",x"fb"),
  3960 => (x"c0",x"1e",x"74",x"87"),
  3961 => (x"87",x"db",x"f9",x"49"),
  3962 => (x"49",x"73",x"1e",x"74"),
  3963 => (x"c8",x"87",x"d4",x"f9"),
  3964 => (x"73",x"87",x"c6",x"86"),
  3965 => (x"cc",x"d0",x"fd",x"49"),
  3966 => (x"87",x"ef",x"fe",x"87"),
  3967 => (x"f9",x"c3",x"1e",x"00"),
  3968 => (x"c1",x"49",x"bf",x"cb"),
  3969 => (x"cf",x"f9",x"c3",x"b9"),
  3970 => (x"48",x"d4",x"ff",x"59"),
  3971 => (x"ff",x"78",x"ff",x"c3"),
  3972 => (x"e1",x"c8",x"48",x"d0"),
  3973 => (x"48",x"d4",x"ff",x"78"),
  3974 => (x"31",x"c4",x"78",x"c1"),
  3975 => (x"d0",x"ff",x"78",x"71"),
  3976 => (x"78",x"e0",x"c0",x"48"),
  3977 => (x"c3",x"1e",x"4f",x"26"),
  3978 => (x"c4",x"1e",x"ff",x"f8"),
  3979 => (x"fc",x"49",x"e6",x"f2"),
  3980 => (x"c4",x"87",x"db",x"ef"),
  3981 => (x"02",x"98",x"70",x"86"),
  3982 => (x"c0",x"ff",x"87",x"c3"),
  3983 => (x"31",x"4f",x"26",x"87"),
  3984 => (x"5a",x"48",x"4b",x"35"),
  3985 => (x"43",x"20",x"20",x"20"),
  3986 => (x"00",x"00",x"47",x"46"),
  3987 => (x"1a",x"00",x"00",x"00"),
  3988 => (x"11",x"12",x"58",x"9f"),
  3989 => (x"1c",x"1b",x"1d",x"14"),
  3990 => (x"5a",x"a7",x"4a",x"23"),
  3991 => (x"f5",x"94",x"91",x"59"),
  3992 => (x"f5",x"f4",x"eb",x"f2"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

