library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"10307c7c",
     1 => x"60301000",
     2 => x"061e7860",
     3 => x"3c664200",
     4 => x"42663c18",
     5 => x"6a387800",
     6 => x"386cc6c2",
     7 => x"00006000",
     8 => x"60000060",
     9 => x"5b5e0e00",
    10 => x"1e0e5d5c",
    11 => x"f0c24c71",
    12 => x"c04dbfc6",
    13 => x"741ec04b",
    14 => x"87c702ab",
    15 => x"c048a6c4",
    16 => x"c487c578",
    17 => x"78c148a6",
    18 => x"731e66c4",
    19 => x"87dfee49",
    20 => x"e0c086c8",
    21 => x"87efef49",
    22 => x"6a4aa5c4",
    23 => x"87f0f049",
    24 => x"cb87c6f1",
    25 => x"c883c185",
    26 => x"ff04abb7",
    27 => x"262687c7",
    28 => x"264c264d",
    29 => x"1e4f264b",
    30 => x"f0c24a71",
    31 => x"f0c25aca",
    32 => x"78c748ca",
    33 => x"87ddfe49",
    34 => x"731e4f26",
    35 => x"c04a711e",
    36 => x"d303aab7",
    37 => x"d1d0c287",
    38 => x"87c405bf",
    39 => x"87c24bc1",
    40 => x"d0c24bc0",
    41 => x"87c45bd5",
    42 => x"5ad5d0c2",
    43 => x"bfd1d0c2",
    44 => x"c19ac14a",
    45 => x"ec49a2c0",
    46 => x"48fc87e8",
    47 => x"bfd1d0c2",
    48 => x"87effe78",
    49 => x"c44a711e",
    50 => x"49721e66",
    51 => x"2687f5e9",
    52 => x"c21e4f26",
    53 => x"49bfd1d0",
    54 => x"c287c8e6",
    55 => x"e848feef",
    56 => x"efc278bf",
    57 => x"bfec48fa",
    58 => x"feefc278",
    59 => x"cf494abf",
    60 => x"b7ca99ff",
    61 => x"7148722a",
    62 => x"c6f0c2b0",
    63 => x"0e4f2658",
    64 => x"5d5c5b5e",
    65 => x"ff4b710e",
    66 => x"efc287c8",
    67 => x"50c048f9",
    68 => x"f5e54973",
    69 => x"4c497087",
    70 => x"eecb9cc2",
    71 => x"87f9cb49",
    72 => x"c24d4970",
    73 => x"bf97f9ef",
    74 => x"87e2c105",
    75 => x"c24966d0",
    76 => x"99bfc2f0",
    77 => x"d487d605",
    78 => x"efc24966",
    79 => x"0599bffa",
    80 => x"497387cb",
    81 => x"7087c3e5",
    82 => x"c1c10298",
    83 => x"fe4cc187",
    84 => x"497587c0",
    85 => x"7087cecb",
    86 => x"87c60298",
    87 => x"48f9efc2",
    88 => x"efc250c1",
    89 => x"05bf97f9",
    90 => x"c287e3c0",
    91 => x"49bfc2f0",
    92 => x"059966d0",
    93 => x"c287d6ff",
    94 => x"49bffaef",
    95 => x"059966d4",
    96 => x"7387caff",
    97 => x"87c2e449",
    98 => x"fe059870",
    99 => x"487487ff",
   100 => x"0e87dcfb",
   101 => x"5d5c5b5e",
   102 => x"c086f40e",
   103 => x"bfec4c4d",
   104 => x"48a6c47e",
   105 => x"bfc6f0c2",
   106 => x"c01ec178",
   107 => x"fd49c71e",
   108 => x"86c887cd",
   109 => x"cd029870",
   110 => x"fb49ff87",
   111 => x"dac187cc",
   112 => x"87c6e349",
   113 => x"efc24dc1",
   114 => x"02bf97f9",
   115 => x"ded587c3",
   116 => x"feefc287",
   117 => x"d0c24bbf",
   118 => x"c105bfd1",
   119 => x"a6c487da",
   120 => x"c0c0c248",
   121 => x"dec278c0",
   122 => x"976e7ec1",
   123 => x"486e49bf",
   124 => x"7e7080c1",
   125 => x"87d2e271",
   126 => x"c3029870",
   127 => x"b366c487",
   128 => x"c14866c4",
   129 => x"a6c828b7",
   130 => x"05987058",
   131 => x"c387dbff",
   132 => x"f5e149fd",
   133 => x"49fac387",
   134 => x"7387efe1",
   135 => x"99ffcf49",
   136 => x"49c01e71",
   137 => x"7387ddfa",
   138 => x"29b7ca49",
   139 => x"49c11e71",
   140 => x"c887d1fa",
   141 => x"87ffc586",
   142 => x"bfc2f0c2",
   143 => x"dd029b4b",
   144 => x"cdd0c287",
   145 => x"dcc749bf",
   146 => x"05987087",
   147 => x"4bc087c4",
   148 => x"e0c287d2",
   149 => x"87c1c749",
   150 => x"58d1d0c2",
   151 => x"d0c287c6",
   152 => x"78c048cd",
   153 => x"99c24973",
   154 => x"c387cd05",
   155 => x"d9e049eb",
   156 => x"c2497087",
   157 => x"87c20299",
   158 => x"49734cfb",
   159 => x"cd0599c1",
   160 => x"49f4c387",
   161 => x"7087c3e0",
   162 => x"0299c249",
   163 => x"4cfa87c2",
   164 => x"99c84973",
   165 => x"c387ce05",
   166 => x"dfff49f5",
   167 => x"497087ec",
   168 => x"d50299c2",
   169 => x"caf0c287",
   170 => x"87ca02bf",
   171 => x"c288c148",
   172 => x"c058cef0",
   173 => x"4cff87c2",
   174 => x"49734dc1",
   175 => x"ce0599c4",
   176 => x"49f2c387",
   177 => x"87c2dfff",
   178 => x"99c24970",
   179 => x"c287dc02",
   180 => x"7ebfcaf0",
   181 => x"a8b7c748",
   182 => x"87cbc003",
   183 => x"80c1486e",
   184 => x"58cef0c2",
   185 => x"fe87c2c0",
   186 => x"c34dc14c",
   187 => x"deff49fd",
   188 => x"497087d8",
   189 => x"c00299c2",
   190 => x"f0c287d5",
   191 => x"c002bfca",
   192 => x"f0c287c9",
   193 => x"78c048ca",
   194 => x"fd87c2c0",
   195 => x"c34dc14c",
   196 => x"ddff49fa",
   197 => x"497087f4",
   198 => x"c00299c2",
   199 => x"f0c287d9",
   200 => x"c748bfca",
   201 => x"c003a8b7",
   202 => x"f0c287c9",
   203 => x"78c748ca",
   204 => x"fc87c2c0",
   205 => x"c04dc14c",
   206 => x"c003acb7",
   207 => x"66c487d1",
   208 => x"82d8c14a",
   209 => x"c6c0026a",
   210 => x"744b6a87",
   211 => x"c00f7349",
   212 => x"1ef0c31e",
   213 => x"f649dac1",
   214 => x"86c887e5",
   215 => x"c0029870",
   216 => x"a6c887e2",
   217 => x"caf0c248",
   218 => x"66c878bf",
   219 => x"c491cb49",
   220 => x"80714866",
   221 => x"bf6e7e70",
   222 => x"87c8c002",
   223 => x"c84bbf6e",
   224 => x"0f734966",
   225 => x"c0029d75",
   226 => x"f0c287c8",
   227 => x"f249bfca",
   228 => x"d0c287d3",
   229 => x"c002bfd5",
   230 => x"c24987dd",
   231 => x"987087c7",
   232 => x"87d3c002",
   233 => x"bfcaf0c2",
   234 => x"87f9f149",
   235 => x"d9f349c0",
   236 => x"d5d0c287",
   237 => x"f478c048",
   238 => x"87f3f28e",
   239 => x"5c5b5e0e",
   240 => x"711e0e5d",
   241 => x"c6f0c24c",
   242 => x"cdc149bf",
   243 => x"d1c14da1",
   244 => x"747e6981",
   245 => x"87cf029c",
   246 => x"744ba5c4",
   247 => x"c6f0c27b",
   248 => x"d2f249bf",
   249 => x"747b6e87",
   250 => x"87c4059c",
   251 => x"87c24bc0",
   252 => x"49734bc1",
   253 => x"d487d3f2",
   254 => x"87c70266",
   255 => x"7087da49",
   256 => x"c087c24a",
   257 => x"d9d0c24a",
   258 => x"e2f1265a",
   259 => x"00000087",
   260 => x"00000000",
   261 => x"00000000",
   262 => x"4a711e00",
   263 => x"49bfc8ff",
   264 => x"2648a172",
   265 => x"c8ff1e4f",
   266 => x"c0fe89bf",
   267 => x"c0c0c0c0",
   268 => x"87c401a9",
   269 => x"87c24ac0",
   270 => x"48724ac1",
   271 => x"5e0e4f26",
   272 => x"0e5d5c5b",
   273 => x"d4ff4b71",
   274 => x"4866d04c",
   275 => x"49d678c0",
   276 => x"87f6daff",
   277 => x"6c7cffc3",
   278 => x"99ffc349",
   279 => x"c3494d71",
   280 => x"e0c199f0",
   281 => x"87cb05a9",
   282 => x"6c7cffc3",
   283 => x"d098c348",
   284 => x"c3780866",
   285 => x"4a6c7cff",
   286 => x"c331c849",
   287 => x"4a6c7cff",
   288 => x"4972b271",
   289 => x"ffc331c8",
   290 => x"714a6c7c",
   291 => x"c84972b2",
   292 => x"7cffc331",
   293 => x"b2714a6c",
   294 => x"c048d0ff",
   295 => x"9b7378e0",
   296 => x"7287c202",
   297 => x"2648757b",
   298 => x"264c264d",
   299 => x"1e4f264b",
   300 => x"5e0e4f26",
   301 => x"f80e5c5b",
   302 => x"c81e7686",
   303 => x"fdfd49a6",
   304 => x"7086c487",
   305 => x"c0486e4b",
   306 => x"f0c201a8",
   307 => x"c34a7387",
   308 => x"d0c19af0",
   309 => x"87c702aa",
   310 => x"05aae0c1",
   311 => x"7387dec2",
   312 => x"0299c849",
   313 => x"c6ff87c3",
   314 => x"c34c7387",
   315 => x"05acc29c",
   316 => x"c487c2c1",
   317 => x"31c94966",
   318 => x"66c41e71",
   319 => x"c292d44a",
   320 => x"7249cef0",
   321 => x"e6d2fe81",
   322 => x"ff49d887",
   323 => x"c887fbd7",
   324 => x"dec21ec0",
   325 => x"effd49fe",
   326 => x"d0ff87c1",
   327 => x"78e0c048",
   328 => x"1efedec2",
   329 => x"d44a66cc",
   330 => x"cef0c292",
   331 => x"fe817249",
   332 => x"cc87f9d0",
   333 => x"05acc186",
   334 => x"c487c2c1",
   335 => x"31c94966",
   336 => x"66c41e71",
   337 => x"c292d44a",
   338 => x"7249cef0",
   339 => x"ded1fe81",
   340 => x"fedec287",
   341 => x"4a66c81e",
   342 => x"f0c292d4",
   343 => x"817249ce",
   344 => x"87c5cffe",
   345 => x"d6ff49d7",
   346 => x"c0c887e0",
   347 => x"fedec21e",
   348 => x"d0edfd49",
   349 => x"ff86cc87",
   350 => x"e0c048d0",
   351 => x"fc8ef878",
   352 => x"5e0e87e7",
   353 => x"0e5d5c5b",
   354 => x"ff4d711e",
   355 => x"66d44cd4",
   356 => x"b7c3487e",
   357 => x"87c506a8",
   358 => x"e2c148c0",
   359 => x"fe497587",
   360 => x"7587dddf",
   361 => x"4b66c41e",
   362 => x"f0c293d4",
   363 => x"497383ce",
   364 => x"87d9cafe",
   365 => x"4b6b83c8",
   366 => x"c848d0ff",
   367 => x"7cdd78e1",
   368 => x"ffc34973",
   369 => x"737c7199",
   370 => x"29b7c849",
   371 => x"7199ffc3",
   372 => x"d049737c",
   373 => x"ffc329b7",
   374 => x"737c7199",
   375 => x"29b7d849",
   376 => x"7cc07c71",
   377 => x"7c7c7c7c",
   378 => x"7c7c7c7c",
   379 => x"c07c7c7c",
   380 => x"66c478e0",
   381 => x"ff49dc1e",
   382 => x"c887f4d4",
   383 => x"26487386",
   384 => x"0e87e4fa",
   385 => x"5d5c5b5e",
   386 => x"7e711e0e",
   387 => x"6e4bd4ff",
   388 => x"e2f0c21e",
   389 => x"f4c8fe49",
   390 => x"7086c487",
   391 => x"c3029d4d",
   392 => x"f0c287c3",
   393 => x"6e4cbfea",
   394 => x"d3ddfe49",
   395 => x"48d0ff87",
   396 => x"c178c5c8",
   397 => x"4ac07bd6",
   398 => x"82c17b15",
   399 => x"aab7e0c0",
   400 => x"ff87f504",
   401 => x"78c448d0",
   402 => x"c178c5c8",
   403 => x"7bc17bd3",
   404 => x"9c7478c4",
   405 => x"87fcc102",
   406 => x"7efedec2",
   407 => x"8c4dc0c8",
   408 => x"03acb7c0",
   409 => x"c0c887c6",
   410 => x"4cc04da4",
   411 => x"97efebc2",
   412 => x"99d049bf",
   413 => x"c087d202",
   414 => x"e2f0c21e",
   415 => x"e8cafe49",
   416 => x"7086c487",
   417 => x"efc04a49",
   418 => x"fedec287",
   419 => x"e2f0c21e",
   420 => x"d4cafe49",
   421 => x"7086c487",
   422 => x"d0ff4a49",
   423 => x"78c5c848",
   424 => x"6e7bd4c1",
   425 => x"6e7bbf97",
   426 => x"7080c148",
   427 => x"058dc17e",
   428 => x"ff87f0ff",
   429 => x"78c448d0",
   430 => x"c5059a72",
   431 => x"c048c087",
   432 => x"1ec187e5",
   433 => x"49e2f0c2",
   434 => x"87fcc7fe",
   435 => x"9c7486c4",
   436 => x"87c4fe05",
   437 => x"c848d0ff",
   438 => x"d3c178c5",
   439 => x"c47bc07b",
   440 => x"c248c178",
   441 => x"2648c087",
   442 => x"4c264d26",
   443 => x"4f264b26",
   444 => x"5c5b5e0e",
   445 => x"cc4b710e",
   446 => x"87d80266",
   447 => x"8cf0c04c",
   448 => x"7487d802",
   449 => x"028ac14a",
   450 => x"028a87d1",
   451 => x"028a87cd",
   452 => x"87d787c9",
   453 => x"eafb4973",
   454 => x"7487d087",
   455 => x"f949c01e",
   456 => x"1e7487e0",
   457 => x"d9f94973",
   458 => x"fe86c887",
   459 => x"1e0087fc",
   460 => x"bffdddc2",
   461 => x"c2b9c149",
   462 => x"ff59c1de",
   463 => x"ffc348d4",
   464 => x"48d0ff78",
   465 => x"ff78e1c8",
   466 => x"78c148d4",
   467 => x"787131c4",
   468 => x"c048d0ff",
   469 => x"4f2678e0",
   470 => x"f1ddc21e",
   471 => x"e2f0c21e",
   472 => x"e8c3fe49",
   473 => x"7086c487",
   474 => x"87c30298",
   475 => x"2687c0ff",
   476 => x"4b35314f",
   477 => x"20205a48",
   478 => x"47464320",
   479 => x"00000000",
   480 => x"589f1a00",
   481 => x"1d141112",
   482 => x"4a231c1b",
   483 => x"91595aa7",
   484 => x"ebf2f594",
   485 => x"ebf2f5f4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
