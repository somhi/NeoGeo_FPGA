library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ecf2c487",
    12 => x"86c0c64e",
    13 => x"49ecf2c4",
    14 => x"48d4f9c3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e3eb",
    19 => x"1e87fc98",
    20 => x"48121e72",
    21 => x"87c40211",
    22 => x"87f60288",
    23 => x"4f264a26",
    24 => x"731e721e",
    25 => x"1148121e",
    26 => x"4b87ca02",
    27 => x"9b98dfc3",
    28 => x"f0028873",
    29 => x"264b2687",
    30 => x"1e4f264a",
    31 => x"1e721e73",
    32 => x"ca048bc1",
    33 => x"11481287",
    34 => x"8887c402",
    35 => x"2687f102",
    36 => x"264b264a",
    37 => x"1e741e4f",
    38 => x"1e721e73",
    39 => x"d0048bc1",
    40 => x"11481287",
    41 => x"4c87ca02",
    42 => x"9c98dfc3",
    43 => x"eb028874",
    44 => x"264a2687",
    45 => x"264c264b",
    46 => x"48731e4f",
    47 => x"02a97381",
    48 => x"531287c5",
    49 => x"2687f605",
    50 => x"66c41e4f",
    51 => x"1248714a",
    52 => x"87fb0551",
    53 => x"731e4f26",
    54 => x"a9738148",
    55 => x"f9537205",
    56 => x"0e4f2687",
    57 => x"5d5c5b5e",
    58 => x"7186f40e",
    59 => x"48a6c44d",
    60 => x"66dc78c0",
    61 => x"48a6c84b",
    62 => x"971578c0",
    63 => x"026e977e",
    64 => x"1387f0c0",
    65 => x"da029c4c",
    66 => x"4a6e9787",
    67 => x"aab74974",
    68 => x"c887c905",
    69 => x"78c148a6",
    70 => x"87c24cc0",
    71 => x"9c744c13",
    72 => x"c887e605",
    73 => x"87cb0266",
    74 => x"c14866c4",
    75 => x"58a6c880",
    76 => x"c487fffe",
    77 => x"8ef44866",
    78 => x"4c264d26",
    79 => x"4f264b26",
    80 => x"c14a711e",
    81 => x"04aab7c1",
    82 => x"c6c187d9",
    83 => x"d201aab7",
    84 => x"4866c487",
    85 => x"ca05a8d0",
    86 => x"c0497287",
    87 => x"487189f7",
    88 => x"c187ecc0",
    89 => x"04aab7e1",
    90 => x"e6c187d8",
    91 => x"d101aab7",
    92 => x"4866c487",
    93 => x"c905a8d0",
    94 => x"c1497287",
    95 => x"487189d7",
    96 => x"f0c087cd",
    97 => x"aab7c98a",
    98 => x"ff87c206",
    99 => x"2648724a",
   100 => x"5b5e0e4f",
   101 => x"f80e5d5c",
   102 => x"c47e7186",
   103 => x"78c048a6",
   104 => x"a7f9c14c",
   105 => x"4966c41e",
   106 => x"c487f8fc",
   107 => x"6e497086",
   108 => x"9783714b",
   109 => x"edc0496b",
   110 => x"87c605a9",
   111 => x"c148a6c4",
   112 => x"66d88378",
   113 => x"d887c502",
   114 => x"0b7b0b66",
   115 => x"d3056b97",
   116 => x"0266c487",
   117 => x"4a7487c7",
   118 => x"c28a0ac0",
   119 => x"724a7487",
   120 => x"87efc048",
   121 => x"131e66dc",
   122 => x"87d4fd49",
   123 => x"4d7086c4",
   124 => x"03adb7c0",
   125 => x"66c487d4",
   126 => x"7487c902",
   127 => x"8808c048",
   128 => x"87c27e70",
   129 => x"486e7e74",
   130 => x"66dc87c9",
   131 => x"4ca47594",
   132 => x"f887effe",
   133 => x"264d268e",
   134 => x"264b264c",
   135 => x"1e00204f",
   136 => x"9a721e73",
   137 => x"87e7c002",
   138 => x"4bc148c0",
   139 => x"d106a972",
   140 => x"06827287",
   141 => x"837387c9",
   142 => x"f401a972",
   143 => x"c187c387",
   144 => x"a9723ab2",
   145 => x"80738903",
   146 => x"2b2ac107",
   147 => x"2687f305",
   148 => x"1e4f264b",
   149 => x"4dc41e75",
   150 => x"04a1b771",
   151 => x"81c1b9ff",
   152 => x"7207bdc3",
   153 => x"ff04a2b7",
   154 => x"c182c1ba",
   155 => x"eefe07bd",
   156 => x"042dc187",
   157 => x"80c1b8ff",
   158 => x"ff042d07",
   159 => x"0781c1b9",
   160 => x"4f264d26",
   161 => x"ff48111e",
   162 => x"c47808d4",
   163 => x"88c14866",
   164 => x"7058a6c8",
   165 => x"87ed0598",
   166 => x"ff1e4f26",
   167 => x"ffc348d4",
   168 => x"c4516878",
   169 => x"88c14866",
   170 => x"7058a6c8",
   171 => x"87eb0598",
   172 => x"731e4f26",
   173 => x"4bd4ff1e",
   174 => x"6b7bffc3",
   175 => x"7bffc34a",
   176 => x"32c8496b",
   177 => x"ffc3b172",
   178 => x"c84a6b7b",
   179 => x"c3b27131",
   180 => x"496b7bff",
   181 => x"b17232c8",
   182 => x"87c44871",
   183 => x"4c264d26",
   184 => x"4f264b26",
   185 => x"5c5b5e0e",
   186 => x"4a710e5d",
   187 => x"724cd4ff",
   188 => x"99ffc349",
   189 => x"f9c37c71",
   190 => x"c805bfd4",
   191 => x"4866d087",
   192 => x"a6d430c9",
   193 => x"4966d058",
   194 => x"ffc329d8",
   195 => x"d07c7199",
   196 => x"29d04966",
   197 => x"7199ffc3",
   198 => x"4966d07c",
   199 => x"ffc329c8",
   200 => x"d07c7199",
   201 => x"ffc34966",
   202 => x"727c7199",
   203 => x"c329d049",
   204 => x"7c7199ff",
   205 => x"f0c94b6c",
   206 => x"ffc34dff",
   207 => x"87d005ab",
   208 => x"6c7cffc3",
   209 => x"028dc14b",
   210 => x"ffc387c6",
   211 => x"87f002ab",
   212 => x"c7fe4873",
   213 => x"49c01e87",
   214 => x"c348d4ff",
   215 => x"81c178ff",
   216 => x"a9b7c8c3",
   217 => x"2687f104",
   218 => x"1e731e4f",
   219 => x"f8c487e7",
   220 => x"1ec04bdf",
   221 => x"c1f0ffc0",
   222 => x"e7fd49f7",
   223 => x"c186c487",
   224 => x"eac005a8",
   225 => x"48d4ff87",
   226 => x"c178ffc3",
   227 => x"c0c0c0c0",
   228 => x"e1c01ec0",
   229 => x"49e9c1f0",
   230 => x"c487c9fd",
   231 => x"05987086",
   232 => x"d4ff87ca",
   233 => x"78ffc348",
   234 => x"87cb48c1",
   235 => x"c187e6fe",
   236 => x"fdfe058b",
   237 => x"fc48c087",
   238 => x"731e87e6",
   239 => x"48d4ff1e",
   240 => x"d378ffc3",
   241 => x"c01ec04b",
   242 => x"c1c1f0ff",
   243 => x"87d4fc49",
   244 => x"987086c4",
   245 => x"ff87ca05",
   246 => x"ffc348d4",
   247 => x"cb48c178",
   248 => x"87f1fd87",
   249 => x"ff058bc1",
   250 => x"48c087db",
   251 => x"0e87f1fb",
   252 => x"0e5c5b5e",
   253 => x"fd4cd4ff",
   254 => x"eac687db",
   255 => x"f0e1c01e",
   256 => x"fb49c8c1",
   257 => x"86c487de",
   258 => x"c802a8c1",
   259 => x"87eafe87",
   260 => x"e2c148c0",
   261 => x"87dafa87",
   262 => x"ffcf4970",
   263 => x"eac699ff",
   264 => x"87c802a9",
   265 => x"c087d3fe",
   266 => x"87cbc148",
   267 => x"c07cffc3",
   268 => x"f4fc4bf1",
   269 => x"02987087",
   270 => x"c087ebc0",
   271 => x"f0ffc01e",
   272 => x"fa49fac1",
   273 => x"86c487de",
   274 => x"d9059870",
   275 => x"7cffc387",
   276 => x"ffc3496c",
   277 => x"7c7c7c7c",
   278 => x"0299c0c1",
   279 => x"48c187c4",
   280 => x"48c087d5",
   281 => x"abc287d1",
   282 => x"c087c405",
   283 => x"c187c848",
   284 => x"fdfe058b",
   285 => x"f948c087",
   286 => x"731e87e4",
   287 => x"d4f9c31e",
   288 => x"c778c148",
   289 => x"48d0ff4b",
   290 => x"c8fb78c2",
   291 => x"48d0ff87",
   292 => x"1ec078c3",
   293 => x"c1d0e5c0",
   294 => x"c7f949c0",
   295 => x"c186c487",
   296 => x"87c105a8",
   297 => x"05abc24b",
   298 => x"48c087c5",
   299 => x"c187f9c0",
   300 => x"d0ff058b",
   301 => x"87f7fc87",
   302 => x"58d8f9c3",
   303 => x"cd059870",
   304 => x"c01ec187",
   305 => x"d0c1f0ff",
   306 => x"87d8f849",
   307 => x"d4ff86c4",
   308 => x"78ffc348",
   309 => x"c387e0c4",
   310 => x"ff58dcf9",
   311 => x"78c248d0",
   312 => x"c348d4ff",
   313 => x"48c178ff",
   314 => x"0e87f5f7",
   315 => x"5d5c5b5e",
   316 => x"c34a710e",
   317 => x"d4ff4dff",
   318 => x"ff7c754c",
   319 => x"c3c448d0",
   320 => x"727c7578",
   321 => x"f0ffc01e",
   322 => x"f749d8c1",
   323 => x"86c487d6",
   324 => x"c5029870",
   325 => x"c048c087",
   326 => x"7c7587f0",
   327 => x"c87cfec3",
   328 => x"66d41ec0",
   329 => x"87dcf549",
   330 => x"7c7586c4",
   331 => x"7c757c75",
   332 => x"4be0dad8",
   333 => x"496c7c75",
   334 => x"87c50599",
   335 => x"f3058bc1",
   336 => x"ff7c7587",
   337 => x"78c248d0",
   338 => x"cff648c1",
   339 => x"d4ff1e87",
   340 => x"48d0ff4a",
   341 => x"c378d1c4",
   342 => x"89c17aff",
   343 => x"2687f805",
   344 => x"1e731e4f",
   345 => x"eec54b71",
   346 => x"ff4adfcd",
   347 => x"ffc348d4",
   348 => x"c3486878",
   349 => x"c502a8fe",
   350 => x"058ac187",
   351 => x"9a7287ed",
   352 => x"c087c505",
   353 => x"87eac048",
   354 => x"cc029b73",
   355 => x"1e66c887",
   356 => x"c5f44973",
   357 => x"c686c487",
   358 => x"4966c887",
   359 => x"ff87eefe",
   360 => x"ffc348d4",
   361 => x"9b737878",
   362 => x"ff87c505",
   363 => x"78d048d0",
   364 => x"ebf448c1",
   365 => x"1e731e87",
   366 => x"4bc04a71",
   367 => x"c348d4ff",
   368 => x"d0ff78ff",
   369 => x"78c3c448",
   370 => x"c348d4ff",
   371 => x"1e7278ff",
   372 => x"c1f0ffc0",
   373 => x"cbf449d1",
   374 => x"7086c487",
   375 => x"87cd0598",
   376 => x"cc1ec0c8",
   377 => x"f8fd4966",
   378 => x"7086c487",
   379 => x"48d0ff4b",
   380 => x"487378c2",
   381 => x"0e87e9f3",
   382 => x"5d5c5b5e",
   383 => x"c01ec00e",
   384 => x"c9c1f0ff",
   385 => x"87dcf349",
   386 => x"f9c31ed2",
   387 => x"d0fd49dc",
   388 => x"c086c887",
   389 => x"d284c14c",
   390 => x"f804acb7",
   391 => x"dcf9c387",
   392 => x"c349bf97",
   393 => x"c0c199c0",
   394 => x"e7c005a9",
   395 => x"e3f9c387",
   396 => x"d049bf97",
   397 => x"e4f9c331",
   398 => x"c84abf97",
   399 => x"c3b17232",
   400 => x"bf97e5f9",
   401 => x"4c71b14a",
   402 => x"ffffffcf",
   403 => x"ca84c19c",
   404 => x"87e7c134",
   405 => x"97e5f9c3",
   406 => x"31c149bf",
   407 => x"f9c399c6",
   408 => x"4abf97e6",
   409 => x"722ab7c7",
   410 => x"e1f9c3b1",
   411 => x"4d4abf97",
   412 => x"f9c39dcf",
   413 => x"4abf97e2",
   414 => x"32ca9ac3",
   415 => x"97e3f9c3",
   416 => x"33c24bbf",
   417 => x"f9c3b273",
   418 => x"4bbf97e4",
   419 => x"c69bc0c3",
   420 => x"b2732bb7",
   421 => x"48c181c2",
   422 => x"49703071",
   423 => x"307548c1",
   424 => x"4c724d70",
   425 => x"947184c1",
   426 => x"adb7c0c8",
   427 => x"c187cc06",
   428 => x"c82db734",
   429 => x"01adb7c0",
   430 => x"7487f4ff",
   431 => x"87dcf048",
   432 => x"5c5b5e0e",
   433 => x"86f80e5d",
   434 => x"48c2c2c4",
   435 => x"f9c378c0",
   436 => x"49c01efa",
   437 => x"c487defb",
   438 => x"05987086",
   439 => x"48c087c5",
   440 => x"c087cec9",
   441 => x"c07ec14d",
   442 => x"49bff9fe",
   443 => x"4af0fac3",
   444 => x"e64bc871",
   445 => x"987087c5",
   446 => x"c087c205",
   447 => x"f5fec07e",
   448 => x"fbc349bf",
   449 => x"c8714acc",
   450 => x"87efe54b",
   451 => x"c2059870",
   452 => x"6e7ec087",
   453 => x"87fdc002",
   454 => x"bfc0c1c4",
   455 => x"f8c1c44d",
   456 => x"487ebf9f",
   457 => x"a8ead6c5",
   458 => x"c487c705",
   459 => x"4dbfc0c1",
   460 => x"486e87ce",
   461 => x"a8d5e9ca",
   462 => x"c087c502",
   463 => x"87f1c748",
   464 => x"1efaf9c3",
   465 => x"ecf94975",
   466 => x"7086c487",
   467 => x"87c50598",
   468 => x"dcc748c0",
   469 => x"f5fec087",
   470 => x"fbc349bf",
   471 => x"c8714acc",
   472 => x"87d7e44b",
   473 => x"c8059870",
   474 => x"c2c2c487",
   475 => x"da78c148",
   476 => x"f9fec087",
   477 => x"fac349bf",
   478 => x"c8714af0",
   479 => x"87fbe34b",
   480 => x"c0029870",
   481 => x"48c087c5",
   482 => x"c487e6c6",
   483 => x"bf97f8c1",
   484 => x"a9d5c149",
   485 => x"87cdc005",
   486 => x"97f9c1c4",
   487 => x"eac249bf",
   488 => x"c5c002a9",
   489 => x"c648c087",
   490 => x"f9c387c7",
   491 => x"7ebf97fa",
   492 => x"a8e9c348",
   493 => x"87cec002",
   494 => x"ebc3486e",
   495 => x"c5c002a8",
   496 => x"c548c087",
   497 => x"fac387eb",
   498 => x"49bf97c5",
   499 => x"ccc00599",
   500 => x"c6fac387",
   501 => x"c249bf97",
   502 => x"c5c002a9",
   503 => x"c548c087",
   504 => x"fac387cf",
   505 => x"48bf97c7",
   506 => x"58fec1c4",
   507 => x"c1484c70",
   508 => x"c2c2c488",
   509 => x"c8fac358",
   510 => x"7549bf97",
   511 => x"c9fac381",
   512 => x"c84abf97",
   513 => x"7ea17232",
   514 => x"48cfc6c4",
   515 => x"fac3786e",
   516 => x"48bf97ca",
   517 => x"c458a6c8",
   518 => x"02bfc2c2",
   519 => x"c087d4c2",
   520 => x"49bff5fe",
   521 => x"4accfbc3",
   522 => x"e14bc871",
   523 => x"987087cd",
   524 => x"87c5c002",
   525 => x"f8c348c0",
   526 => x"fac1c487",
   527 => x"c6c44cbf",
   528 => x"fac35ce3",
   529 => x"49bf97df",
   530 => x"fac331c8",
   531 => x"4abf97de",
   532 => x"fac349a1",
   533 => x"4abf97e0",
   534 => x"a17232d0",
   535 => x"e1fac349",
   536 => x"d84abf97",
   537 => x"49a17232",
   538 => x"c49166c4",
   539 => x"81bfcfc6",
   540 => x"59d7c6c4",
   541 => x"97e7fac3",
   542 => x"32c84abf",
   543 => x"97e6fac3",
   544 => x"4aa24bbf",
   545 => x"97e8fac3",
   546 => x"33d04bbf",
   547 => x"c34aa273",
   548 => x"bf97e9fa",
   549 => x"d89bcf4b",
   550 => x"4aa27333",
   551 => x"5adbc6c4",
   552 => x"bfd7c6c4",
   553 => x"748ac24a",
   554 => x"dbc6c492",
   555 => x"78a17248",
   556 => x"c387cac1",
   557 => x"bf97ccfa",
   558 => x"c331c849",
   559 => x"bf97cbfa",
   560 => x"c449a14a",
   561 => x"c459cac2",
   562 => x"49bfc6c2",
   563 => x"ffc731c5",
   564 => x"c429c981",
   565 => x"c359e3c6",
   566 => x"bf97d1fa",
   567 => x"c332c84a",
   568 => x"bf97d0fa",
   569 => x"c44aa24b",
   570 => x"826e9266",
   571 => x"5adfc6c4",
   572 => x"48d7c6c4",
   573 => x"c6c478c0",
   574 => x"a17248d3",
   575 => x"e3c6c478",
   576 => x"d7c6c448",
   577 => x"c6c478bf",
   578 => x"c6c448e7",
   579 => x"c478bfdb",
   580 => x"02bfc2c2",
   581 => x"7487c9c0",
   582 => x"7030c448",
   583 => x"87c9c07e",
   584 => x"bfdfc6c4",
   585 => x"7030c448",
   586 => x"c6c2c47e",
   587 => x"c1786e48",
   588 => x"268ef848",
   589 => x"264c264d",
   590 => x"0e4f264b",
   591 => x"5d5c5b5e",
   592 => x"c44a710e",
   593 => x"02bfc2c2",
   594 => x"4b7287cb",
   595 => x"4c722bc7",
   596 => x"c99cffc1",
   597 => x"c84b7287",
   598 => x"c34c722b",
   599 => x"c6c49cff",
   600 => x"c083bfcf",
   601 => x"abbff1fe",
   602 => x"c087d902",
   603 => x"c35bf5fe",
   604 => x"731efaf9",
   605 => x"87fdf049",
   606 => x"987086c4",
   607 => x"c087c505",
   608 => x"87e6c048",
   609 => x"bfc2c2c4",
   610 => x"7487d202",
   611 => x"c391c449",
   612 => x"6981faf9",
   613 => x"ffffcf4d",
   614 => x"cb9dffff",
   615 => x"c2497487",
   616 => x"faf9c391",
   617 => x"4d699f81",
   618 => x"c6fe4875",
   619 => x"5b5e0e87",
   620 => x"1e0e5d5c",
   621 => x"1ec04d71",
   622 => x"dcd049c1",
   623 => x"7086c487",
   624 => x"c1029c4c",
   625 => x"c2c487c2",
   626 => x"49754aca",
   627 => x"87d0daff",
   628 => x"c0029870",
   629 => x"4a7487f2",
   630 => x"4bcb4975",
   631 => x"87f5daff",
   632 => x"c0029870",
   633 => x"1ec087e2",
   634 => x"c7029c74",
   635 => x"48a6c487",
   636 => x"87c578c0",
   637 => x"c148a6c4",
   638 => x"4966c478",
   639 => x"c487dacf",
   640 => x"9c4c7086",
   641 => x"87fefe05",
   642 => x"fc264874",
   643 => x"5e0e87e5",
   644 => x"0e5d5c5b",
   645 => x"9b4b711e",
   646 => x"c087c505",
   647 => x"87e5c148",
   648 => x"c04da3c8",
   649 => x"0266d47d",
   650 => x"66d487c7",
   651 => x"c505bf97",
   652 => x"c148c087",
   653 => x"66d487cf",
   654 => x"87f1fd49",
   655 => x"029c4c70",
   656 => x"dc87c0c1",
   657 => x"7d6949a4",
   658 => x"c449a4da",
   659 => x"699f4aa3",
   660 => x"c2c2c47a",
   661 => x"87d202bf",
   662 => x"9f49a4d4",
   663 => x"ffc04969",
   664 => x"487199ff",
   665 => x"7e7030d0",
   666 => x"7ec087c2",
   667 => x"6a48496e",
   668 => x"c07a7080",
   669 => x"49a3cc7b",
   670 => x"a3d0796a",
   671 => x"7479c049",
   672 => x"c087c248",
   673 => x"eafa2648",
   674 => x"5b5e0e87",
   675 => x"710e5d5c",
   676 => x"f1fec04c",
   677 => x"7478ff48",
   678 => x"cac1029c",
   679 => x"49a4c887",
   680 => x"c2c10269",
   681 => x"4a66d087",
   682 => x"d482496c",
   683 => x"66d05aa6",
   684 => x"c1c4b94d",
   685 => x"ff4abffe",
   686 => x"719972ba",
   687 => x"e4c00299",
   688 => x"4ba4c487",
   689 => x"f2f9496b",
   690 => x"c47b7087",
   691 => x"49bffac1",
   692 => x"7c71816c",
   693 => x"c1c4b975",
   694 => x"ff4abffe",
   695 => x"719972ba",
   696 => x"dcff0599",
   697 => x"f97c7587",
   698 => x"731e87c9",
   699 => x"9b4b711e",
   700 => x"c887c702",
   701 => x"056949a3",
   702 => x"48c087c5",
   703 => x"c487ebc0",
   704 => x"4abfd3c6",
   705 => x"6949a3c4",
   706 => x"c489c249",
   707 => x"91bffac1",
   708 => x"c44aa271",
   709 => x"49bffec1",
   710 => x"a271996b",
   711 => x"1e66c84a",
   712 => x"d0ea4972",
   713 => x"7086c487",
   714 => x"caf84849",
   715 => x"1e731e87",
   716 => x"029b4b71",
   717 => x"a3c887c7",
   718 => x"c5056949",
   719 => x"c048c087",
   720 => x"c6c487eb",
   721 => x"c44abfd3",
   722 => x"496949a3",
   723 => x"c1c489c2",
   724 => x"7191bffa",
   725 => x"c1c44aa2",
   726 => x"6b49bffe",
   727 => x"4aa27199",
   728 => x"721e66c8",
   729 => x"87c3e649",
   730 => x"497086c4",
   731 => x"87c7f748",
   732 => x"5c5b5e0e",
   733 => x"711e0e5d",
   734 => x"4c66d44b",
   735 => x"9b732cc9",
   736 => x"87cfc102",
   737 => x"6949a3c8",
   738 => x"87c7c102",
   739 => x"d44da3d0",
   740 => x"c1c47d66",
   741 => x"ff49bffe",
   742 => x"994a6bb9",
   743 => x"03ac717e",
   744 => x"7bc087cd",
   745 => x"4aa3cc7d",
   746 => x"6a49a3c4",
   747 => x"7287c279",
   748 => x"029c748c",
   749 => x"1e4987dd",
   750 => x"ccfb4973",
   751 => x"d486c487",
   752 => x"ffc74966",
   753 => x"87cb0299",
   754 => x"1efaf9c3",
   755 => x"d9fc4973",
   756 => x"2686c487",
   757 => x"0e87dcf5",
   758 => x"5d5c5b5e",
   759 => x"d086f00e",
   760 => x"e4c059a6",
   761 => x"66cc4b66",
   762 => x"4887ca02",
   763 => x"7e7080c8",
   764 => x"c505bf6e",
   765 => x"c348c087",
   766 => x"66cc87ec",
   767 => x"7384d04c",
   768 => x"48a6c449",
   769 => x"66c4786c",
   770 => x"6e80c481",
   771 => x"66c878bf",
   772 => x"87c606a9",
   773 => x"8966c449",
   774 => x"b7c04b71",
   775 => x"87c401ab",
   776 => x"87c2c348",
   777 => x"c74866c4",
   778 => x"7e7098ff",
   779 => x"c9c1026e",
   780 => x"49c0c887",
   781 => x"4a71896e",
   782 => x"4dfaf9c3",
   783 => x"b773856e",
   784 => x"87c106aa",
   785 => x"4849724a",
   786 => x"708066c4",
   787 => x"498b727c",
   788 => x"99718ac1",
   789 => x"c087d902",
   790 => x"154866e0",
   791 => x"66e0c050",
   792 => x"c080c148",
   793 => x"7258a6e4",
   794 => x"718ac149",
   795 => x"87e70599",
   796 => x"66d01ec1",
   797 => x"87d1f849",
   798 => x"b7c086c4",
   799 => x"e3c106ab",
   800 => x"66e0c087",
   801 => x"b7ffc74d",
   802 => x"e2c006ab",
   803 => x"d01e7587",
   804 => x"d5f94966",
   805 => x"85c0c887",
   806 => x"c0c8486c",
   807 => x"c87c7080",
   808 => x"1ec18bc0",
   809 => x"f74966d4",
   810 => x"86c887df",
   811 => x"c387eec0",
   812 => x"d01efaf9",
   813 => x"f1f84966",
   814 => x"c386c487",
   815 => x"734afaf9",
   816 => x"806c4849",
   817 => x"49737c70",
   818 => x"99718bc1",
   819 => x"1287ce02",
   820 => x"85c17d97",
   821 => x"8bc14973",
   822 => x"f2059971",
   823 => x"abb7c087",
   824 => x"87e1fe01",
   825 => x"8ef048c1",
   826 => x"0e87c8f1",
   827 => x"5d5c5b5e",
   828 => x"9b4b710e",
   829 => x"c887c702",
   830 => x"056d4da3",
   831 => x"48ff87c5",
   832 => x"d087fdc0",
   833 => x"496c4ca3",
   834 => x"0599ffc7",
   835 => x"026c87d8",
   836 => x"1ec187c9",
   837 => x"f0f54973",
   838 => x"c386c487",
   839 => x"731efaf9",
   840 => x"87c6f749",
   841 => x"4a6c86c4",
   842 => x"c404aa6d",
   843 => x"cf48ff87",
   844 => x"7ca2c187",
   845 => x"ffc74972",
   846 => x"faf9c399",
   847 => x"48699781",
   848 => x"1e87f0ef",
   849 => x"4b711e73",
   850 => x"e4c0029b",
   851 => x"e7c6c487",
   852 => x"c24a735b",
   853 => x"fac1c48a",
   854 => x"c49249bf",
   855 => x"48bfd3c6",
   856 => x"c6c48072",
   857 => x"487158eb",
   858 => x"c2c430c4",
   859 => x"edc058ca",
   860 => x"e3c6c487",
   861 => x"d7c6c448",
   862 => x"c6c478bf",
   863 => x"c6c448e7",
   864 => x"c478bfdb",
   865 => x"02bfc2c2",
   866 => x"c1c487c9",
   867 => x"c449bffa",
   868 => x"c487c731",
   869 => x"49bfdfc6",
   870 => x"c2c431c4",
   871 => x"d6ee59ca",
   872 => x"5b5e0e87",
   873 => x"4a710e5c",
   874 => x"9a724bc0",
   875 => x"87e1c002",
   876 => x"9f49a2da",
   877 => x"c2c44b69",
   878 => x"cf02bfc2",
   879 => x"49a2d487",
   880 => x"4c49699f",
   881 => x"9cffffc0",
   882 => x"87c234d0",
   883 => x"49744cc0",
   884 => x"fd4973b3",
   885 => x"dced87ed",
   886 => x"5b5e0e87",
   887 => x"f40e5d5c",
   888 => x"c04a7186",
   889 => x"029a727e",
   890 => x"f9c387d8",
   891 => x"78c048f6",
   892 => x"48eef9c3",
   893 => x"bfe7c6c4",
   894 => x"f2f9c378",
   895 => x"e3c6c448",
   896 => x"c2c478bf",
   897 => x"50c048d7",
   898 => x"bfc6c2c4",
   899 => x"f6f9c349",
   900 => x"aa714abf",
   901 => x"87c0c403",
   902 => x"99cf4972",
   903 => x"87e1c005",
   904 => x"1efaf9c3",
   905 => x"bfeef9c3",
   906 => x"eef9c349",
   907 => x"78a1c148",
   908 => x"c0deff71",
   909 => x"c086c487",
   910 => x"c348edfe",
   911 => x"cc78faf9",
   912 => x"edfec087",
   913 => x"e0c048bf",
   914 => x"f1fec080",
   915 => x"f6f9c358",
   916 => x"80c148bf",
   917 => x"58faf9c3",
   918 => x"000fad27",
   919 => x"bf97bf00",
   920 => x"c2029d4d",
   921 => x"e5c387e2",
   922 => x"dbc202ad",
   923 => x"edfec087",
   924 => x"a3cb4bbf",
   925 => x"cf4c1149",
   926 => x"d2c105ac",
   927 => x"df497587",
   928 => x"cd89c199",
   929 => x"cac2c491",
   930 => x"4aa3c181",
   931 => x"a3c35112",
   932 => x"c551124a",
   933 => x"51124aa3",
   934 => x"124aa3c7",
   935 => x"4aa3c951",
   936 => x"a3ce5112",
   937 => x"d051124a",
   938 => x"51124aa3",
   939 => x"124aa3d2",
   940 => x"4aa3d451",
   941 => x"a3d65112",
   942 => x"d851124a",
   943 => x"51124aa3",
   944 => x"124aa3dc",
   945 => x"4aa3de51",
   946 => x"7ec15112",
   947 => x"7487f9c0",
   948 => x"0599c849",
   949 => x"7487eac0",
   950 => x"0599d049",
   951 => x"66dc87d0",
   952 => x"87cac002",
   953 => x"66dc4973",
   954 => x"0298700f",
   955 => x"056e87d3",
   956 => x"c487c6c0",
   957 => x"c048cac2",
   958 => x"edfec050",
   959 => x"e7c248bf",
   960 => x"d7c2c487",
   961 => x"7e50c048",
   962 => x"bfc6c2c4",
   963 => x"f6f9c349",
   964 => x"aa714abf",
   965 => x"87c0fc04",
   966 => x"bfe7c6c4",
   967 => x"87c8c005",
   968 => x"bfc2c2c4",
   969 => x"87fec102",
   970 => x"48f1fec0",
   971 => x"f9c378ff",
   972 => x"e849bff2",
   973 => x"497087c5",
   974 => x"59f6f9c3",
   975 => x"c348a6c4",
   976 => x"78bff2f9",
   977 => x"bfc2c2c4",
   978 => x"87d8c002",
   979 => x"cf4966c4",
   980 => x"f8ffffff",
   981 => x"c002a999",
   982 => x"4dc087c5",
   983 => x"c187e1c0",
   984 => x"87dcc04d",
   985 => x"cf4966c4",
   986 => x"a999f8ff",
   987 => x"87c8c002",
   988 => x"c048a6c8",
   989 => x"87c5c078",
   990 => x"c148a6c8",
   991 => x"4d66c878",
   992 => x"c0059d75",
   993 => x"66c487e0",
   994 => x"c489c249",
   995 => x"4abffac1",
   996 => x"d3c6c491",
   997 => x"f9c34abf",
   998 => x"a17248ee",
   999 => x"f6f9c378",
  1000 => x"f978c048",
  1001 => x"48c087e2",
  1002 => x"c6e68ef4",
  1003 => x"00000087",
  1004 => x"ffffff00",
  1005 => x"000fbdff",
  1006 => x"000fc600",
  1007 => x"54414600",
  1008 => x"20203233",
  1009 => x"41460020",
  1010 => x"20363154",
  1011 => x"1e002020",
  1012 => x"c348d4ff",
  1013 => x"486878ff",
  1014 => x"ff1e4f26",
  1015 => x"ffc348d4",
  1016 => x"48d0ff78",
  1017 => x"ff78e1c8",
  1018 => x"78d448d4",
  1019 => x"48ebc6c4",
  1020 => x"50bfd4ff",
  1021 => x"ff1e4f26",
  1022 => x"e0c048d0",
  1023 => x"1e4f2678",
  1024 => x"7087ccff",
  1025 => x"c6029949",
  1026 => x"a9fbc087",
  1027 => x"7187f105",
  1028 => x"0e4f2648",
  1029 => x"0e5c5b5e",
  1030 => x"4cc04b71",
  1031 => x"7087f0fe",
  1032 => x"c0029949",
  1033 => x"ecc087f9",
  1034 => x"f2c002a9",
  1035 => x"a9fbc087",
  1036 => x"87ebc002",
  1037 => x"acb766cc",
  1038 => x"d087c703",
  1039 => x"87c20266",
  1040 => x"99715371",
  1041 => x"c187c202",
  1042 => x"87c3fe84",
  1043 => x"02994970",
  1044 => x"ecc087cd",
  1045 => x"87c702a9",
  1046 => x"05a9fbc0",
  1047 => x"d087d5ff",
  1048 => x"87c30266",
  1049 => x"c07b97c0",
  1050 => x"c405a9ec",
  1051 => x"c54a7487",
  1052 => x"c04a7487",
  1053 => x"48728a0a",
  1054 => x"4d2687c2",
  1055 => x"4b264c26",
  1056 => x"fd1e4f26",
  1057 => x"497087c9",
  1058 => x"a9b7f0c0",
  1059 => x"c087ca04",
  1060 => x"01a9b7f9",
  1061 => x"f0c087c3",
  1062 => x"b7c1c189",
  1063 => x"87ca04a9",
  1064 => x"a9b7dac1",
  1065 => x"c087c301",
  1066 => x"487189f7",
  1067 => x"5e0e4f26",
  1068 => x"710e5c5b",
  1069 => x"4cd4ff4a",
  1070 => x"eac04972",
  1071 => x"9b4b7087",
  1072 => x"c187c202",
  1073 => x"48d0ff8b",
  1074 => x"c178c5c8",
  1075 => x"49737cd5",
  1076 => x"f7c331c6",
  1077 => x"4abf97eb",
  1078 => x"70b07148",
  1079 => x"48d0ff7c",
  1080 => x"487378c4",
  1081 => x"0e87d5fe",
  1082 => x"5d5c5b5e",
  1083 => x"7186f80e",
  1084 => x"fb7ec04c",
  1085 => x"4bc087e4",
  1086 => x"97d4c6c1",
  1087 => x"a9c049bf",
  1088 => x"fb87cf04",
  1089 => x"83c187f9",
  1090 => x"97d4c6c1",
  1091 => x"06ab49bf",
  1092 => x"c6c187f1",
  1093 => x"02bf97d4",
  1094 => x"f2fa87cf",
  1095 => x"99497087",
  1096 => x"c087c602",
  1097 => x"f105a9ec",
  1098 => x"fa4bc087",
  1099 => x"4d7087e1",
  1100 => x"c887dcfa",
  1101 => x"d6fa58a6",
  1102 => x"c14a7087",
  1103 => x"49a4c883",
  1104 => x"ad496997",
  1105 => x"c087c702",
  1106 => x"c005adff",
  1107 => x"a4c987e7",
  1108 => x"49699749",
  1109 => x"02a966c4",
  1110 => x"c04887c7",
  1111 => x"d405a8ff",
  1112 => x"49a4ca87",
  1113 => x"aa496997",
  1114 => x"c087c602",
  1115 => x"c405aaff",
  1116 => x"d07ec187",
  1117 => x"adecc087",
  1118 => x"c087c602",
  1119 => x"c405adfb",
  1120 => x"c14bc087",
  1121 => x"fe026e7e",
  1122 => x"e9f987e1",
  1123 => x"f8487387",
  1124 => x"87e6fb8e",
  1125 => x"5b5e0e00",
  1126 => x"1e0e5d5c",
  1127 => x"4cc04b71",
  1128 => x"c004ab4d",
  1129 => x"c3c187e8",
  1130 => x"9d751ee7",
  1131 => x"c087c402",
  1132 => x"c187c24a",
  1133 => x"f049724a",
  1134 => x"86c487df",
  1135 => x"84c17e70",
  1136 => x"87c2056e",
  1137 => x"85c14c73",
  1138 => x"ff06ac73",
  1139 => x"486e87d8",
  1140 => x"264d2626",
  1141 => x"264b264c",
  1142 => x"4a711e4f",
  1143 => x"99ffc349",
  1144 => x"7148d4ff",
  1145 => x"c8497278",
  1146 => x"ffc329b7",
  1147 => x"72787199",
  1148 => x"29b7d049",
  1149 => x"7199ffc3",
  1150 => x"d8497278",
  1151 => x"ffc329b7",
  1152 => x"26787199",
  1153 => x"5b5e0e4f",
  1154 => x"1e0e5d5c",
  1155 => x"4bc04a71",
  1156 => x"e3c14972",
  1157 => x"987087c5",
  1158 => x"c187da05",
  1159 => x"c149744c",
  1160 => x"7087d2e4",
  1161 => x"87c20598",
  1162 => x"84c14bc1",
  1163 => x"bfcecbc4",
  1164 => x"e806acb7",
  1165 => x"48d0ff87",
  1166 => x"ff78e1c8",
  1167 => x"78dd48d4",
  1168 => x"c7029b73",
  1169 => x"f6cbc487",
  1170 => x"87c24dbf",
  1171 => x"49754dc0",
  1172 => x"7387c6fe",
  1173 => x"87c7029b",
  1174 => x"bff6cbc4",
  1175 => x"c087c27e",
  1176 => x"fd496e7e",
  1177 => x"49c087f3",
  1178 => x"c087eefd",
  1179 => x"87e9fd49",
  1180 => x"c048d0ff",
  1181 => x"1ec178e0",
  1182 => x"f2c049dc",
  1183 => x"487387ca",
  1184 => x"ccfd8ef8",
  1185 => x"5b5e0e87",
  1186 => x"1e0e5d5c",
  1187 => x"de494c71",
  1188 => x"c5c7c491",
  1189 => x"9785714d",
  1190 => x"ddc1026d",
  1191 => x"f0c6c487",
  1192 => x"82744abf",
  1193 => x"ecfb4972",
  1194 => x"6e7e7087",
  1195 => x"87f3c002",
  1196 => x"4bf8c6c4",
  1197 => x"49cb4a6e",
  1198 => x"87fdf7fe",
  1199 => x"93cb4b74",
  1200 => x"83d3edc1",
  1201 => x"cbc183c4",
  1202 => x"49747bfe",
  1203 => x"87eec4c1",
  1204 => x"c7c47b75",
  1205 => x"49bf97c4",
  1206 => x"f8c6c41e",
  1207 => x"ffeac249",
  1208 => x"7486c487",
  1209 => x"d5c4c149",
  1210 => x"c149c087",
  1211 => x"c487f4c5",
  1212 => x"c048ecc6",
  1213 => x"dd49c178",
  1214 => x"fb2687c1",
  1215 => x"6f4c87d3",
  1216 => x"6e696461",
  1217 => x"2e2e2e67",
  1218 => x"5b5e0e00",
  1219 => x"4b710e5c",
  1220 => x"f0c6c44a",
  1221 => x"497282bf",
  1222 => x"7087faf9",
  1223 => x"c4029c4c",
  1224 => x"fce94987",
  1225 => x"f0c6c487",
  1226 => x"c178c048",
  1227 => x"87cbdc49",
  1228 => x"0e87e0fa",
  1229 => x"5d5c5b5e",
  1230 => x"c386f40e",
  1231 => x"c04dfaf9",
  1232 => x"48a6c44c",
  1233 => x"c6c478c0",
  1234 => x"c049bff0",
  1235 => x"c1c106a9",
  1236 => x"faf9c387",
  1237 => x"c0029848",
  1238 => x"c3c187f8",
  1239 => x"66c81ee7",
  1240 => x"c487c702",
  1241 => x"78c048a6",
  1242 => x"a6c487c5",
  1243 => x"c478c148",
  1244 => x"e4e94966",
  1245 => x"7086c487",
  1246 => x"c484c14d",
  1247 => x"80c14866",
  1248 => x"c458a6c8",
  1249 => x"49bff0c6",
  1250 => x"87c603ac",
  1251 => x"ff059d75",
  1252 => x"4cc087c8",
  1253 => x"c3029d75",
  1254 => x"c3c187e0",
  1255 => x"66c81ee7",
  1256 => x"cc87c702",
  1257 => x"78c048a6",
  1258 => x"a6cc87c5",
  1259 => x"cc78c148",
  1260 => x"e4e84966",
  1261 => x"7086c487",
  1262 => x"c2026e7e",
  1263 => x"496e87e9",
  1264 => x"699781cb",
  1265 => x"0299d049",
  1266 => x"c187d6c1",
  1267 => x"744ac9cc",
  1268 => x"c191cb49",
  1269 => x"7281d3ed",
  1270 => x"c381c879",
  1271 => x"497451ff",
  1272 => x"c7c491de",
  1273 => x"85714dc5",
  1274 => x"7d97c1c2",
  1275 => x"c049a5c1",
  1276 => x"c2c451e0",
  1277 => x"02bf97ca",
  1278 => x"84c187d2",
  1279 => x"c44ba5c2",
  1280 => x"db4acac2",
  1281 => x"f0f2fe49",
  1282 => x"87dbc187",
  1283 => x"c049a5cd",
  1284 => x"c284c151",
  1285 => x"4a6e4ba5",
  1286 => x"f2fe49cb",
  1287 => x"c6c187db",
  1288 => x"c5cac187",
  1289 => x"cb49744a",
  1290 => x"d3edc191",
  1291 => x"c4797281",
  1292 => x"bf97cac2",
  1293 => x"7487d802",
  1294 => x"c191de49",
  1295 => x"c5c7c484",
  1296 => x"c483714b",
  1297 => x"dd4acac2",
  1298 => x"ecf1fe49",
  1299 => x"7487d887",
  1300 => x"c493de4b",
  1301 => x"cb83c5c7",
  1302 => x"51c049a3",
  1303 => x"6e7384c1",
  1304 => x"fe49cb4a",
  1305 => x"c487d2f1",
  1306 => x"80c14866",
  1307 => x"c758a6c8",
  1308 => x"c5c003ac",
  1309 => x"fc056e87",
  1310 => x"487487e0",
  1311 => x"d0f58ef4",
  1312 => x"1e731e87",
  1313 => x"cb494b71",
  1314 => x"d3edc191",
  1315 => x"4aa1c881",
  1316 => x"48ebf7c3",
  1317 => x"a1c95012",
  1318 => x"d4c6c14a",
  1319 => x"ca501248",
  1320 => x"c4c7c481",
  1321 => x"c4501148",
  1322 => x"bf97c4c7",
  1323 => x"49c01e49",
  1324 => x"87ece3c2",
  1325 => x"48ecc6c4",
  1326 => x"49c178de",
  1327 => x"2687fcd5",
  1328 => x"1e87d2f4",
  1329 => x"cb494a71",
  1330 => x"d3edc191",
  1331 => x"1181c881",
  1332 => x"f0c6c448",
  1333 => x"f0c6c458",
  1334 => x"c178c048",
  1335 => x"87dbd549",
  1336 => x"c01e4f26",
  1337 => x"fafdc049",
  1338 => x"1e4f2687",
  1339 => x"d2029971",
  1340 => x"e8eec187",
  1341 => x"f750c048",
  1342 => x"c3d3c180",
  1343 => x"ccedc140",
  1344 => x"c187ce78",
  1345 => x"c148e4ee",
  1346 => x"fc78c5ed",
  1347 => x"e2d3c180",
  1348 => x"0e4f2678",
  1349 => x"0e5c5b5e",
  1350 => x"cb4a4c71",
  1351 => x"d3edc192",
  1352 => x"49a2c882",
  1353 => x"974ba2c9",
  1354 => x"971e4b6b",
  1355 => x"ca1e4969",
  1356 => x"c0491282",
  1357 => x"c087f5e8",
  1358 => x"87ffd349",
  1359 => x"fac04974",
  1360 => x"8ef887fc",
  1361 => x"1e87ccf2",
  1362 => x"4b711e73",
  1363 => x"87c3ff49",
  1364 => x"fefe4973",
  1365 => x"87fdf187",
  1366 => x"711e731e",
  1367 => x"4aa3c64b",
  1368 => x"c187db02",
  1369 => x"87d6028a",
  1370 => x"dac1028a",
  1371 => x"c0028a87",
  1372 => x"028a87fc",
  1373 => x"8a87e1c0",
  1374 => x"c187cb02",
  1375 => x"49c787db",
  1376 => x"c187c0fd",
  1377 => x"c6c487de",
  1378 => x"c102bff0",
  1379 => x"c14887cb",
  1380 => x"f4c6c488",
  1381 => x"87c1c158",
  1382 => x"bff4c6c4",
  1383 => x"87f9c002",
  1384 => x"bff0c6c4",
  1385 => x"c480c148",
  1386 => x"c058f4c6",
  1387 => x"c6c487eb",
  1388 => x"c649bff0",
  1389 => x"f4c6c489",
  1390 => x"a9b7c059",
  1391 => x"c487da03",
  1392 => x"c048f0c6",
  1393 => x"c487d278",
  1394 => x"02bff4c6",
  1395 => x"c6c487cb",
  1396 => x"c648bff0",
  1397 => x"f4c6c480",
  1398 => x"d149c058",
  1399 => x"497387dd",
  1400 => x"87daf8c0",
  1401 => x"0e87eeef",
  1402 => x"0e5c5b5e",
  1403 => x"66cc4c71",
  1404 => x"cb4b741e",
  1405 => x"d3edc193",
  1406 => x"4aa3c483",
  1407 => x"ebfe496a",
  1408 => x"d2c187c7",
  1409 => x"a3c87bc1",
  1410 => x"5166d449",
  1411 => x"d849a3c9",
  1412 => x"a3ca5166",
  1413 => x"5166dc49",
  1414 => x"87f7ee26",
  1415 => x"5c5b5e0e",
  1416 => x"d0ff0e5d",
  1417 => x"59a6d886",
  1418 => x"c048a6c4",
  1419 => x"c180c478",
  1420 => x"c47866c4",
  1421 => x"c478c180",
  1422 => x"c478c180",
  1423 => x"c148f4c6",
  1424 => x"ecc6c478",
  1425 => x"a8de48bf",
  1426 => x"f387cb05",
  1427 => x"497087e5",
  1428 => x"ce59a6c8",
  1429 => x"c1e687ed",
  1430 => x"87e3e687",
  1431 => x"7087f0e5",
  1432 => x"acfbc04c",
  1433 => x"87d0c102",
  1434 => x"c10566d4",
  1435 => x"1ec087c2",
  1436 => x"c11ec11e",
  1437 => x"c01ec6ef",
  1438 => x"87ebfd49",
  1439 => x"4a66d0c1",
  1440 => x"496a82c4",
  1441 => x"517481c7",
  1442 => x"1ed81ec1",
  1443 => x"81c8496a",
  1444 => x"d887c0e6",
  1445 => x"66c4c186",
  1446 => x"01a8c048",
  1447 => x"a6c487c7",
  1448 => x"ce78c148",
  1449 => x"66c4c187",
  1450 => x"cc88c148",
  1451 => x"87c358a6",
  1452 => x"cc87cce5",
  1453 => x"78c248a6",
  1454 => x"cd029c74",
  1455 => x"66c487c1",
  1456 => x"66c8c148",
  1457 => x"f6cc03a8",
  1458 => x"48a6d887",
  1459 => x"80c478c0",
  1460 => x"fae378c0",
  1461 => x"c14c7087",
  1462 => x"c205acd0",
  1463 => x"66dc87d7",
  1464 => x"87dee67e",
  1465 => x"e0c04970",
  1466 => x"e2e359a6",
  1467 => x"c04c7087",
  1468 => x"c105acec",
  1469 => x"66c487ea",
  1470 => x"c191cb49",
  1471 => x"c48166c0",
  1472 => x"4d6a4aa1",
  1473 => x"dc4aa1c8",
  1474 => x"d3c15266",
  1475 => x"fee279c3",
  1476 => x"9c4c7087",
  1477 => x"c087d802",
  1478 => x"d202acfb",
  1479 => x"e2557487",
  1480 => x"4c7087ed",
  1481 => x"87c7029c",
  1482 => x"05acfbc0",
  1483 => x"c087eeff",
  1484 => x"c1c255e0",
  1485 => x"7d97c055",
  1486 => x"6e4966d4",
  1487 => x"87db05a9",
  1488 => x"c84866c4",
  1489 => x"ca04a866",
  1490 => x"4866c487",
  1491 => x"a6c880c1",
  1492 => x"c887c858",
  1493 => x"88c14866",
  1494 => x"e158a6cc",
  1495 => x"4c7087f1",
  1496 => x"05acd0c1",
  1497 => x"66d087c8",
  1498 => x"d480c148",
  1499 => x"d0c158a6",
  1500 => x"e9fd02ac",
  1501 => x"a6e0c087",
  1502 => x"7866d448",
  1503 => x"c04866dc",
  1504 => x"05a866e0",
  1505 => x"c087cac9",
  1506 => x"c048a6e4",
  1507 => x"48747e78",
  1508 => x"c088fbc0",
  1509 => x"7058a6ec",
  1510 => x"cfc80298",
  1511 => x"88cb4887",
  1512 => x"58a6ecc0",
  1513 => x"c1029870",
  1514 => x"c94887d2",
  1515 => x"a6ecc088",
  1516 => x"02987058",
  1517 => x"4887dbc3",
  1518 => x"ecc088c4",
  1519 => x"987058a6",
  1520 => x"4887d002",
  1521 => x"ecc088c1",
  1522 => x"987058a6",
  1523 => x"87c2c302",
  1524 => x"d887d3c7",
  1525 => x"f0c048a6",
  1526 => x"f2dfff78",
  1527 => x"c04c7087",
  1528 => x"c002acec",
  1529 => x"a6dc87c3",
  1530 => x"acecc05c",
  1531 => x"ff87cd02",
  1532 => x"7087dcdf",
  1533 => x"acecc04c",
  1534 => x"87f3ff05",
  1535 => x"02acecc0",
  1536 => x"ff87c4c0",
  1537 => x"d887c8df",
  1538 => x"66d41e66",
  1539 => x"66d41e49",
  1540 => x"efc11e49",
  1541 => x"66d41ec6",
  1542 => x"87cbf749",
  1543 => x"1eca1ec0",
  1544 => x"cb4966dc",
  1545 => x"66d8c191",
  1546 => x"48a6d881",
  1547 => x"d878a1c4",
  1548 => x"ff49bf66",
  1549 => x"d887dcdf",
  1550 => x"a8b7c086",
  1551 => x"87c5c106",
  1552 => x"1ede1ec1",
  1553 => x"49bf66c8",
  1554 => x"87c7dfff",
  1555 => x"497086c8",
  1556 => x"8808c048",
  1557 => x"c058a6dc",
  1558 => x"c006a8b7",
  1559 => x"66d887e7",
  1560 => x"a8b7dd48",
  1561 => x"6e87de03",
  1562 => x"66d849bf",
  1563 => x"51e0c081",
  1564 => x"c14966d8",
  1565 => x"81bf6e81",
  1566 => x"d851c1c2",
  1567 => x"81c24966",
  1568 => x"c081bf6e",
  1569 => x"4866cc51",
  1570 => x"a6d080c1",
  1571 => x"c47ec158",
  1572 => x"dfff87da",
  1573 => x"a6dc87ec",
  1574 => x"e5dfff58",
  1575 => x"a6ecc087",
  1576 => x"a8ecc058",
  1577 => x"87cac005",
  1578 => x"48a6e8c0",
  1579 => x"c07866d8",
  1580 => x"dcff87c4",
  1581 => x"66c487d9",
  1582 => x"c191cb49",
  1583 => x"714866c0",
  1584 => x"6e7e7080",
  1585 => x"6e82c84a",
  1586 => x"d881ca49",
  1587 => x"e8c05166",
  1588 => x"81c14966",
  1589 => x"c18966d8",
  1590 => x"70307148",
  1591 => x"7189c149",
  1592 => x"cac47a97",
  1593 => x"d849bfe1",
  1594 => x"6a972966",
  1595 => x"9871484a",
  1596 => x"58a6f0c0",
  1597 => x"81c4496e",
  1598 => x"e0c04d69",
  1599 => x"66dc4866",
  1600 => x"c8c002a8",
  1601 => x"48a6d887",
  1602 => x"c5c078c0",
  1603 => x"48a6d887",
  1604 => x"66d878c1",
  1605 => x"1ee0c01e",
  1606 => x"dbff4975",
  1607 => x"86c887f5",
  1608 => x"b7c04c70",
  1609 => x"d4c106ac",
  1610 => x"c0857487",
  1611 => x"897449e0",
  1612 => x"e8c14b75",
  1613 => x"fe714af8",
  1614 => x"c287fedd",
  1615 => x"66e4c085",
  1616 => x"c080c148",
  1617 => x"c058a6e8",
  1618 => x"c14966ec",
  1619 => x"02a97081",
  1620 => x"d887c8c0",
  1621 => x"78c048a6",
  1622 => x"d887c5c0",
  1623 => x"78c148a6",
  1624 => x"c21e66d8",
  1625 => x"e0c049a4",
  1626 => x"70887148",
  1627 => x"49751e49",
  1628 => x"87dfdaff",
  1629 => x"b7c086c8",
  1630 => x"c0ff01a8",
  1631 => x"66e4c087",
  1632 => x"87d1c002",
  1633 => x"81c9496e",
  1634 => x"5166e4c0",
  1635 => x"d4c1486e",
  1636 => x"ccc078d3",
  1637 => x"c9496e87",
  1638 => x"6e51c281",
  1639 => x"c7d5c148",
  1640 => x"c07ec178",
  1641 => x"d9ff87c6",
  1642 => x"4c7087d5",
  1643 => x"f5c0026e",
  1644 => x"4866c487",
  1645 => x"04a866c8",
  1646 => x"c487cbc0",
  1647 => x"80c14866",
  1648 => x"c058a6c8",
  1649 => x"66c887e0",
  1650 => x"cc88c148",
  1651 => x"d5c058a6",
  1652 => x"acc6c187",
  1653 => x"87c8c005",
  1654 => x"c14866cc",
  1655 => x"58a6d080",
  1656 => x"87dbd8ff",
  1657 => x"66d04c70",
  1658 => x"d480c148",
  1659 => x"9c7458a6",
  1660 => x"87cbc002",
  1661 => x"c14866c4",
  1662 => x"04a866c8",
  1663 => x"ff87caf3",
  1664 => x"c487f3d7",
  1665 => x"a8c74866",
  1666 => x"87e5c003",
  1667 => x"48f4c6c4",
  1668 => x"66c478c0",
  1669 => x"c191cb49",
  1670 => x"c48166c0",
  1671 => x"4a6a4aa1",
  1672 => x"c47952c0",
  1673 => x"80c14866",
  1674 => x"c758a6c8",
  1675 => x"dbff04a8",
  1676 => x"8ed0ff87",
  1677 => x"87d9deff",
  1678 => x"1e00203a",
  1679 => x"4b711e73",
  1680 => x"87c6029b",
  1681 => x"48f0c6c4",
  1682 => x"1ec778c0",
  1683 => x"bff0c6c4",
  1684 => x"edc11e49",
  1685 => x"c6c41ed3",
  1686 => x"ee49bfec",
  1687 => x"86cc87fe",
  1688 => x"bfecc6c4",
  1689 => x"87c3ea49",
  1690 => x"c8029b73",
  1691 => x"d3edc187",
  1692 => x"dbe7c049",
  1693 => x"dcddff87",
  1694 => x"1e731e87",
  1695 => x"f7c34bc0",
  1696 => x"50c048eb",
  1697 => x"bff6eec1",
  1698 => x"e6c8c249",
  1699 => x"05987087",
  1700 => x"eac187c4",
  1701 => x"48734bdc",
  1702 => x"87f9dcff",
  1703 => x"204d4f52",
  1704 => x"64616f6c",
  1705 => x"20676e69",
  1706 => x"6c696166",
  1707 => x"1e006465",
  1708 => x"c187f2c7",
  1709 => x"87c3fe49",
  1710 => x"87fee6fe",
  1711 => x"cd029870",
  1712 => x"fbeffe87",
  1713 => x"02987087",
  1714 => x"4ac187c4",
  1715 => x"4ac087c2",
  1716 => x"ce059a72",
  1717 => x"c11ec087",
  1718 => x"c049c3ec",
  1719 => x"c487c1f3",
  1720 => x"c287fe86",
  1721 => x"c087eecc",
  1722 => x"ceecc11e",
  1723 => x"eff2c049",
  1724 => x"fe1ec087",
  1725 => x"497087c3",
  1726 => x"87e4f2c0",
  1727 => x"f887e5c3",
  1728 => x"534f268e",
  1729 => x"61662044",
  1730 => x"64656c69",
  1731 => x"6f42002e",
  1732 => x"6e69746f",
  1733 => x"2e2e2e67",
  1734 => x"fcc11e00",
  1735 => x"e9c087c2",
  1736 => x"fbc187cc",
  1737 => x"c0c287fa",
  1738 => x"87ee87f8",
  1739 => x"c41e4f26",
  1740 => x"c048f0c6",
  1741 => x"ecc6c478",
  1742 => x"fd78c048",
  1743 => x"d8ff87f1",
  1744 => x"2648c087",
  1745 => x"4520804f",
  1746 => x"00746978",
  1747 => x"61422080",
  1748 => x"c3006b63",
  1749 => x"c5000014",
  1750 => x"00000041",
  1751 => x"14c30000",
  1752 => x"41e30000",
  1753 => x"00000000",
  1754 => x"0014c300",
  1755 => x"00420100",
  1756 => x"00000000",
  1757 => x"000014c3",
  1758 => x"0000421f",
  1759 => x"c3000000",
  1760 => x"3d000014",
  1761 => x"00000042",
  1762 => x"14c30000",
  1763 => x"425b0000",
  1764 => x"00000000",
  1765 => x"0014c300",
  1766 => x"00427900",
  1767 => x"00000000",
  1768 => x"000014c3",
  1769 => x"00000000",
  1770 => x"58000000",
  1771 => x"00000015",
  1772 => x"00000000",
  1773 => x"1bba0000",
  1774 => x"454e0000",
  1775 => x"4f45474f",
  1776 => x"4f522020",
  1777 => x"6f4c004d",
  1778 => x"2a206461",
  1779 => x"fe1e002e",
  1780 => x"78c048f0",
  1781 => x"097909cd",
  1782 => x"1e1e4f26",
  1783 => x"7ebff0fe",
  1784 => x"4f262648",
  1785 => x"48f0fe1e",
  1786 => x"4f2678c1",
  1787 => x"48f0fe1e",
  1788 => x"4f2678c0",
  1789 => x"c04a711e",
  1790 => x"4f265252",
  1791 => x"5c5b5e0e",
  1792 => x"86f40e5d",
  1793 => x"6d974d71",
  1794 => x"4ca5c17e",
  1795 => x"c8486c97",
  1796 => x"486e58a6",
  1797 => x"05a866c4",
  1798 => x"48ff87c5",
  1799 => x"ff87e6c0",
  1800 => x"a5c287ca",
  1801 => x"4b6c9749",
  1802 => x"974ba371",
  1803 => x"6c974b6b",
  1804 => x"c1486e7e",
  1805 => x"58a6c880",
  1806 => x"a6cc98c7",
  1807 => x"7c977058",
  1808 => x"7387e1fe",
  1809 => x"268ef448",
  1810 => x"264c264d",
  1811 => x"0e4f264b",
  1812 => x"0e5c5b5e",
  1813 => x"4c7186f4",
  1814 => x"c34a66d8",
  1815 => x"a4c29aff",
  1816 => x"496c974b",
  1817 => x"7249a173",
  1818 => x"7e6c9751",
  1819 => x"80c1486e",
  1820 => x"c758a6c8",
  1821 => x"58a6cc98",
  1822 => x"8ef45470",
  1823 => x"1e87caff",
  1824 => x"87e8fd1e",
  1825 => x"494abfe0",
  1826 => x"99c0e0c0",
  1827 => x"7287cb02",
  1828 => x"d7cac41e",
  1829 => x"87f7fe49",
  1830 => x"fdfc86c4",
  1831 => x"fd7e7087",
  1832 => x"262687c2",
  1833 => x"cac41e4f",
  1834 => x"c7fd49d7",
  1835 => x"fff1c187",
  1836 => x"87dafc49",
  1837 => x"2687d5c6",
  1838 => x"5b5e0e4f",
  1839 => x"c40e5d5c",
  1840 => x"4abff6ca",
  1841 => x"bfcdf4c1",
  1842 => x"bc724c49",
  1843 => x"dbfc4d71",
  1844 => x"744bc087",
  1845 => x"0299d049",
  1846 => x"497587d5",
  1847 => x"1e7199d0",
  1848 => x"fbc11ec0",
  1849 => x"82734adb",
  1850 => x"cac14912",
  1851 => x"c186c887",
  1852 => x"c8832d2c",
  1853 => x"daff04ab",
  1854 => x"87e8fb87",
  1855 => x"48cdf4c1",
  1856 => x"bff6cac4",
  1857 => x"264d2678",
  1858 => x"264b264c",
  1859 => x"0000004f",
  1860 => x"1e731e00",
  1861 => x"4ac04b71",
  1862 => x"49dbfbc1",
  1863 => x"69978172",
  1864 => x"05a97349",
  1865 => x"48c187c4",
  1866 => x"82c187ca",
  1867 => x"04aab7c8",
  1868 => x"48c087e6",
  1869 => x"1e87d2ff",
  1870 => x"4b711e73",
  1871 => x"87d1ff49",
  1872 => x"c0029870",
  1873 => x"d0ff87ec",
  1874 => x"78e1c848",
  1875 => x"c548d4ff",
  1876 => x"0266c878",
  1877 => x"e0c387c3",
  1878 => x"0266cc78",
  1879 => x"d4ff87c6",
  1880 => x"78f0c348",
  1881 => x"7348d4ff",
  1882 => x"48d0ff78",
  1883 => x"c078e1c8",
  1884 => x"d4fe78e0",
  1885 => x"5b5e0e87",
  1886 => x"4c710e5c",
  1887 => x"49d7cac4",
  1888 => x"7087f9f9",
  1889 => x"aab7c04a",
  1890 => x"87e3c204",
  1891 => x"05aae0c3",
  1892 => x"f8c187c9",
  1893 => x"78c148f8",
  1894 => x"c387d4c2",
  1895 => x"c905aaf0",
  1896 => x"f4f8c187",
  1897 => x"c178c148",
  1898 => x"f8c187f5",
  1899 => x"c702bff8",
  1900 => x"c24b7287",
  1901 => x"87c2b3c0",
  1902 => x"9c744b72",
  1903 => x"c187d105",
  1904 => x"1ebff4f8",
  1905 => x"bff8f8c1",
  1906 => x"fd49721e",
  1907 => x"86c887e9",
  1908 => x"bff4f8c1",
  1909 => x"87e0c002",
  1910 => x"b7c44973",
  1911 => x"fac19129",
  1912 => x"4a7381db",
  1913 => x"92c29acf",
  1914 => x"307248c1",
  1915 => x"baff4a70",
  1916 => x"98694872",
  1917 => x"87db7970",
  1918 => x"b7c44973",
  1919 => x"fac19129",
  1920 => x"4a7381db",
  1921 => x"92c29acf",
  1922 => x"307248c3",
  1923 => x"69484a70",
  1924 => x"c17970b0",
  1925 => x"c048f8f8",
  1926 => x"f4f8c178",
  1927 => x"c478c048",
  1928 => x"f749d7ca",
  1929 => x"4a7087d6",
  1930 => x"03aab7c0",
  1931 => x"c087ddfd",
  1932 => x"87d3fb48",
  1933 => x"00000000",
  1934 => x"00000000",
  1935 => x"711e731e",
  1936 => x"87f5f94b",
  1937 => x"ecfc4973",
  1938 => x"87fdfa87",
  1939 => x"724ac01e",
  1940 => x"c191c449",
  1941 => x"c081dbfa",
  1942 => x"d082c179",
  1943 => x"ee04aab7",
  1944 => x"0e4f2687",
  1945 => x"5d5c5b5e",
  1946 => x"f54d710e",
  1947 => x"4a7587fe",
  1948 => x"922ab7c4",
  1949 => x"82dbfac1",
  1950 => x"9ccf4c75",
  1951 => x"496a94c2",
  1952 => x"c32b744b",
  1953 => x"7448c29b",
  1954 => x"ff4c7030",
  1955 => x"714874bc",
  1956 => x"f57a7098",
  1957 => x"487387ce",
  1958 => x"0087eaf9",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"16000000",
  1975 => x"2e25261e",
  1976 => x"1e3e3d36",
  1977 => x"c848d0ff",
  1978 => x"487178e1",
  1979 => x"7808d4ff",
  1980 => x"ff1e4f26",
  1981 => x"e1c848d0",
  1982 => x"ff487178",
  1983 => x"c47808d4",
  1984 => x"d4ff4866",
  1985 => x"4f267808",
  1986 => x"c44a711e",
  1987 => x"721e4966",
  1988 => x"87deff49",
  1989 => x"c048d0ff",
  1990 => x"262678e0",
  1991 => x"4a711e4f",
  1992 => x"c11e66c4",
  1993 => x"ff49a2e0",
  1994 => x"66c887c8",
  1995 => x"29b7c849",
  1996 => x"7148d4ff",
  1997 => x"48d0ff78",
  1998 => x"2678e0c0",
  1999 => x"ff1e4f26",
  2000 => x"ffc34ad4",
  2001 => x"48d0ff7a",
  2002 => x"de78e1c8",
  2003 => x"e1cac47a",
  2004 => x"48497abf",
  2005 => x"7a7028c8",
  2006 => x"28d04871",
  2007 => x"48717a70",
  2008 => x"7a7028d8",
  2009 => x"c048d0ff",
  2010 => x"4f2678e0",
  2011 => x"5c5b5e0e",
  2012 => x"4c710e5d",
  2013 => x"bfe1cac4",
  2014 => x"2b744b4d",
  2015 => x"c19b66d0",
  2016 => x"ab66d483",
  2017 => x"c087c204",
  2018 => x"d04a744b",
  2019 => x"31724966",
  2020 => x"9975b9ff",
  2021 => x"30724873",
  2022 => x"71484a70",
  2023 => x"e5cac4b0",
  2024 => x"87dafe58",
  2025 => x"4c264d26",
  2026 => x"4f264b26",
  2027 => x"48d0ff1e",
  2028 => x"7178c9c8",
  2029 => x"08d4ff48",
  2030 => x"1e4f2678",
  2031 => x"eb494a71",
  2032 => x"48d0ff87",
  2033 => x"4f2678c8",
  2034 => x"711e731e",
  2035 => x"f1cac44b",
  2036 => x"87c302bf",
  2037 => x"ff87ebc2",
  2038 => x"c9c848d0",
  2039 => x"c0497378",
  2040 => x"d4ffb1e0",
  2041 => x"c4787148",
  2042 => x"c048e5ca",
  2043 => x"0266c878",
  2044 => x"ffc387c5",
  2045 => x"c087c249",
  2046 => x"edcac449",
  2047 => x"0266cc59",
  2048 => x"d5c587c6",
  2049 => x"87c44ad5",
  2050 => x"4affffcf",
  2051 => x"5af1cac4",
  2052 => x"48f1cac4",
  2053 => x"87c478c1",
  2054 => x"4c264d26",
  2055 => x"4f264b26",
  2056 => x"5c5b5e0e",
  2057 => x"4a710e5d",
  2058 => x"bfedcac4",
  2059 => x"029a724c",
  2060 => x"c84987cb",
  2061 => x"fefec191",
  2062 => x"c483714b",
  2063 => x"fec2c287",
  2064 => x"134dc04b",
  2065 => x"c4997449",
  2066 => x"b9bfe9ca",
  2067 => x"7148d4ff",
  2068 => x"2cb7c178",
  2069 => x"adb7c885",
  2070 => x"c487e804",
  2071 => x"48bfe5ca",
  2072 => x"cac480c8",
  2073 => x"effe58e9",
  2074 => x"1e731e87",
  2075 => x"4a134b71",
  2076 => x"87cb029a",
  2077 => x"e7fe4972",
  2078 => x"9a4a1387",
  2079 => x"fe87f505",
  2080 => x"c41e87da",
  2081 => x"49bfe5ca",
  2082 => x"48e5cac4",
  2083 => x"c478a1c1",
  2084 => x"03a9b7c0",
  2085 => x"d4ff87db",
  2086 => x"e9cac448",
  2087 => x"cac478bf",
  2088 => x"c449bfe5",
  2089 => x"c148e5ca",
  2090 => x"c0c478a1",
  2091 => x"e504a9b7",
  2092 => x"48d0ff87",
  2093 => x"cac478c8",
  2094 => x"78c048f1",
  2095 => x"00004f26",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"005f5f00",
  2099 => x"03000000",
  2100 => x"03030003",
  2101 => x"7f140000",
  2102 => x"7f7f147f",
  2103 => x"24000014",
  2104 => x"3a6b6b2e",
  2105 => x"6a4c0012",
  2106 => x"566c1836",
  2107 => x"7e300032",
  2108 => x"3a77594f",
  2109 => x"00004068",
  2110 => x"00030704",
  2111 => x"00000000",
  2112 => x"41633e1c",
  2113 => x"00000000",
  2114 => x"1c3e6341",
  2115 => x"2a080000",
  2116 => x"3e1c1c3e",
  2117 => x"0800082a",
  2118 => x"083e3e08",
  2119 => x"00000008",
  2120 => x"0060e080",
  2121 => x"08000000",
  2122 => x"08080808",
  2123 => x"00000008",
  2124 => x"00606000",
  2125 => x"60400000",
  2126 => x"060c1830",
  2127 => x"3e000103",
  2128 => x"7f4d597f",
  2129 => x"0400003e",
  2130 => x"007f7f06",
  2131 => x"42000000",
  2132 => x"4f597163",
  2133 => x"22000046",
  2134 => x"7f494963",
  2135 => x"1c180036",
  2136 => x"7f7f1316",
  2137 => x"27000010",
  2138 => x"7d454567",
  2139 => x"3c000039",
  2140 => x"79494b7e",
  2141 => x"01000030",
  2142 => x"0f797101",
  2143 => x"36000007",
  2144 => x"7f49497f",
  2145 => x"06000036",
  2146 => x"3f69494f",
  2147 => x"0000001e",
  2148 => x"00666600",
  2149 => x"00000000",
  2150 => x"0066e680",
  2151 => x"08000000",
  2152 => x"22141408",
  2153 => x"14000022",
  2154 => x"14141414",
  2155 => x"22000014",
  2156 => x"08141422",
  2157 => x"02000008",
  2158 => x"0f595103",
  2159 => x"7f3e0006",
  2160 => x"1f555d41",
  2161 => x"7e00001e",
  2162 => x"7f09097f",
  2163 => x"7f00007e",
  2164 => x"7f49497f",
  2165 => x"1c000036",
  2166 => x"4141633e",
  2167 => x"7f000041",
  2168 => x"3e63417f",
  2169 => x"7f00001c",
  2170 => x"4149497f",
  2171 => x"7f000041",
  2172 => x"0109097f",
  2173 => x"3e000001",
  2174 => x"7b49417f",
  2175 => x"7f00007a",
  2176 => x"7f08087f",
  2177 => x"0000007f",
  2178 => x"417f7f41",
  2179 => x"20000000",
  2180 => x"7f404060",
  2181 => x"7f7f003f",
  2182 => x"63361c08",
  2183 => x"7f000041",
  2184 => x"4040407f",
  2185 => x"7f7f0040",
  2186 => x"7f060c06",
  2187 => x"7f7f007f",
  2188 => x"7f180c06",
  2189 => x"3e00007f",
  2190 => x"7f41417f",
  2191 => x"7f00003e",
  2192 => x"0f09097f",
  2193 => x"7f3e0006",
  2194 => x"7e7f6141",
  2195 => x"7f000040",
  2196 => x"7f19097f",
  2197 => x"26000066",
  2198 => x"7b594d6f",
  2199 => x"01000032",
  2200 => x"017f7f01",
  2201 => x"3f000001",
  2202 => x"7f40407f",
  2203 => x"0f00003f",
  2204 => x"3f70703f",
  2205 => x"7f7f000f",
  2206 => x"7f301830",
  2207 => x"6341007f",
  2208 => x"361c1c36",
  2209 => x"03014163",
  2210 => x"067c7c06",
  2211 => x"71610103",
  2212 => x"43474d59",
  2213 => x"00000041",
  2214 => x"41417f7f",
  2215 => x"03010000",
  2216 => x"30180c06",
  2217 => x"00004060",
  2218 => x"7f7f4141",
  2219 => x"0c080000",
  2220 => x"0c060306",
  2221 => x"80800008",
  2222 => x"80808080",
  2223 => x"00000080",
  2224 => x"04070300",
  2225 => x"20000000",
  2226 => x"7c545474",
  2227 => x"7f000078",
  2228 => x"7c44447f",
  2229 => x"38000038",
  2230 => x"4444447c",
  2231 => x"38000000",
  2232 => x"7f44447c",
  2233 => x"3800007f",
  2234 => x"5c54547c",
  2235 => x"04000018",
  2236 => x"05057f7e",
  2237 => x"18000000",
  2238 => x"fca4a4bc",
  2239 => x"7f00007c",
  2240 => x"7c04047f",
  2241 => x"00000078",
  2242 => x"407d3d00",
  2243 => x"80000000",
  2244 => x"7dfd8080",
  2245 => x"7f000000",
  2246 => x"6c38107f",
  2247 => x"00000044",
  2248 => x"407f3f00",
  2249 => x"7c7c0000",
  2250 => x"7c0c180c",
  2251 => x"7c000078",
  2252 => x"7c04047c",
  2253 => x"38000078",
  2254 => x"7c44447c",
  2255 => x"fc000038",
  2256 => x"3c2424fc",
  2257 => x"18000018",
  2258 => x"fc24243c",
  2259 => x"7c0000fc",
  2260 => x"0c04047c",
  2261 => x"48000008",
  2262 => x"7454545c",
  2263 => x"04000020",
  2264 => x"44447f3f",
  2265 => x"3c000000",
  2266 => x"7c40407c",
  2267 => x"1c00007c",
  2268 => x"3c60603c",
  2269 => x"7c3c001c",
  2270 => x"7c603060",
  2271 => x"6c44003c",
  2272 => x"6c381038",
  2273 => x"1c000044",
  2274 => x"3c60e0bc",
  2275 => x"4400001c",
  2276 => x"4c5c7464",
  2277 => x"08000044",
  2278 => x"41773e08",
  2279 => x"00000041",
  2280 => x"007f7f00",
  2281 => x"41000000",
  2282 => x"083e7741",
  2283 => x"01020008",
  2284 => x"02020301",
  2285 => x"7f7f0001",
  2286 => x"7f7f7f7f",
  2287 => x"0808007f",
  2288 => x"3e3e1c1c",
  2289 => x"7f7f7f7f",
  2290 => x"1c1c3e3e",
  2291 => x"10000808",
  2292 => x"187c7c18",
  2293 => x"10000010",
  2294 => x"307c7c30",
  2295 => x"30100010",
  2296 => x"1e786060",
  2297 => x"66420006",
  2298 => x"663c183c",
  2299 => x"38780042",
  2300 => x"6cc6c26a",
  2301 => x"00600038",
  2302 => x"00006000",
  2303 => x"5e0e0060",
  2304 => x"0e5d5c5b",
  2305 => x"c44c711e",
  2306 => x"4dbfc2cb",
  2307 => x"1ec04bc0",
  2308 => x"c702ab74",
  2309 => x"48a6c487",
  2310 => x"87c578c0",
  2311 => x"c148a6c4",
  2312 => x"1e66c478",
  2313 => x"dfee4973",
  2314 => x"c086c887",
  2315 => x"efef49e0",
  2316 => x"4aa5c487",
  2317 => x"f0f0496a",
  2318 => x"87c6f187",
  2319 => x"83c185cb",
  2320 => x"04abb7c8",
  2321 => x"2687c7ff",
  2322 => x"4c264d26",
  2323 => x"4f264b26",
  2324 => x"c44a711e",
  2325 => x"c45ac6cb",
  2326 => x"c748c6cb",
  2327 => x"ddfe4978",
  2328 => x"1e4f2687",
  2329 => x"4a711e73",
  2330 => x"03aab7c0",
  2331 => x"dfc287d3",
  2332 => x"c405bff7",
  2333 => x"c24bc187",
  2334 => x"c24bc087",
  2335 => x"c45bfbdf",
  2336 => x"fbdfc287",
  2337 => x"f7dfc25a",
  2338 => x"9ac14abf",
  2339 => x"49a2c0c1",
  2340 => x"fc87e8ec",
  2341 => x"f7dfc248",
  2342 => x"effe78bf",
  2343 => x"4a711e87",
  2344 => x"721e66c4",
  2345 => x"87f5e949",
  2346 => x"1e4f2626",
  2347 => x"bff7dfc2",
  2348 => x"87c8e649",
  2349 => x"48facac4",
  2350 => x"c478bfe8",
  2351 => x"ec48f6ca",
  2352 => x"cac478bf",
  2353 => x"494abffa",
  2354 => x"ca99ffcf",
  2355 => x"48722ab7",
  2356 => x"cbc4b071",
  2357 => x"4f2658c2",
  2358 => x"5c5b5e0e",
  2359 => x"4b710e5d",
  2360 => x"c487c8ff",
  2361 => x"c048f5ca",
  2362 => x"e5497350",
  2363 => x"497087f5",
  2364 => x"cb9cc24c",
  2365 => x"d7c149ee",
  2366 => x"497087cf",
  2367 => x"f5cac44d",
  2368 => x"c105bf97",
  2369 => x"66d087e3",
  2370 => x"fecac449",
  2371 => x"d60599bf",
  2372 => x"4966d487",
  2373 => x"bff6cac4",
  2374 => x"87cb0599",
  2375 => x"c2e54973",
  2376 => x"02987087",
  2377 => x"c187c2c1",
  2378 => x"87fffd4c",
  2379 => x"d6c14975",
  2380 => x"987087e3",
  2381 => x"c487c602",
  2382 => x"c148f5ca",
  2383 => x"f5cac450",
  2384 => x"c005bf97",
  2385 => x"cac487e3",
  2386 => x"d049bffe",
  2387 => x"ff059966",
  2388 => x"cac487d5",
  2389 => x"d449bff6",
  2390 => x"ff059966",
  2391 => x"497387c9",
  2392 => x"7087c0e4",
  2393 => x"fefe0598",
  2394 => x"fb487487",
  2395 => x"5e0e87da",
  2396 => x"0e5d5c5b",
  2397 => x"4dc086f4",
  2398 => x"7ebfec4c",
  2399 => x"c448a6c4",
  2400 => x"78bfc2cb",
  2401 => x"1ec01ec1",
  2402 => x"cbfd49c7",
  2403 => x"7086c887",
  2404 => x"87cd0298",
  2405 => x"cafb49ff",
  2406 => x"49dac187",
  2407 => x"c187c4e3",
  2408 => x"f5cac44d",
  2409 => x"c402bf97",
  2410 => x"ffe0c187",
  2411 => x"facac487",
  2412 => x"dfc24bbf",
  2413 => x"c105bff7",
  2414 => x"a6c487da",
  2415 => x"c0c0c248",
  2416 => x"f8c378c0",
  2417 => x"976e7efe",
  2418 => x"486e49bf",
  2419 => x"7e7080c1",
  2420 => x"87cfe271",
  2421 => x"c3029870",
  2422 => x"b366c487",
  2423 => x"c14866c4",
  2424 => x"a6c828b7",
  2425 => x"05987058",
  2426 => x"c387dbff",
  2427 => x"f2e149fd",
  2428 => x"49fac387",
  2429 => x"7387ece1",
  2430 => x"99ffcf49",
  2431 => x"49c01e71",
  2432 => x"7387dafa",
  2433 => x"29b7ca49",
  2434 => x"49c11e71",
  2435 => x"c887cefa",
  2436 => x"87c7c686",
  2437 => x"bffecac4",
  2438 => x"df029b4b",
  2439 => x"f3dfc287",
  2440 => x"d2c149bf",
  2441 => x"987087ef",
  2442 => x"c087c405",
  2443 => x"c287d34b",
  2444 => x"d2c149e0",
  2445 => x"dfc287d3",
  2446 => x"87c658f7",
  2447 => x"48f3dfc2",
  2448 => x"497378c0",
  2449 => x"ce0599c2",
  2450 => x"49ebc387",
  2451 => x"7087d4e0",
  2452 => x"0299c249",
  2453 => x"fb87c2c0",
  2454 => x"c149734c",
  2455 => x"87cf0599",
  2456 => x"ff49f4c3",
  2457 => x"7087fcdf",
  2458 => x"0299c249",
  2459 => x"fa87c2c0",
  2460 => x"c849734c",
  2461 => x"87ce0599",
  2462 => x"ff49f5c3",
  2463 => x"7087e4df",
  2464 => x"0299c249",
  2465 => x"cbc487d6",
  2466 => x"c002bfc6",
  2467 => x"c14887ca",
  2468 => x"cacbc488",
  2469 => x"87c2c058",
  2470 => x"4dc14cff",
  2471 => x"99c44973",
  2472 => x"87cec005",
  2473 => x"ff49f2c3",
  2474 => x"7087f8de",
  2475 => x"0299c249",
  2476 => x"cbc487dc",
  2477 => x"487ebfc6",
  2478 => x"03a8b7c7",
  2479 => x"6e87cbc0",
  2480 => x"c480c148",
  2481 => x"c058cacb",
  2482 => x"4cfe87c2",
  2483 => x"fdc34dc1",
  2484 => x"cedeff49",
  2485 => x"c2497087",
  2486 => x"d5c00299",
  2487 => x"c6cbc487",
  2488 => x"c9c002bf",
  2489 => x"c6cbc487",
  2490 => x"c078c048",
  2491 => x"4cfd87c2",
  2492 => x"fac34dc1",
  2493 => x"eaddff49",
  2494 => x"c2497087",
  2495 => x"d9c00299",
  2496 => x"c6cbc487",
  2497 => x"b7c748bf",
  2498 => x"c9c003a8",
  2499 => x"c6cbc487",
  2500 => x"c078c748",
  2501 => x"4cfc87c2",
  2502 => x"b7c04dc1",
  2503 => x"d1c003ac",
  2504 => x"4a66c487",
  2505 => x"6a82d8c1",
  2506 => x"87c6c002",
  2507 => x"49744b6a",
  2508 => x"1ec00f73",
  2509 => x"c11ef0c3",
  2510 => x"dbf649da",
  2511 => x"7086c887",
  2512 => x"e2c00298",
  2513 => x"48a6c887",
  2514 => x"bfc6cbc4",
  2515 => x"4966c878",
  2516 => x"66c491cb",
  2517 => x"70807148",
  2518 => x"02bf6e7e",
  2519 => x"6e87c8c0",
  2520 => x"66c84bbf",
  2521 => x"750f7349",
  2522 => x"c8c0029d",
  2523 => x"c6cbc487",
  2524 => x"c9f249bf",
  2525 => x"fbdfc287",
  2526 => x"dec002bf",
  2527 => x"cdc14987",
  2528 => x"987087d3",
  2529 => x"87d3c002",
  2530 => x"bfc6cbc4",
  2531 => x"87eef149",
  2532 => x"cef349c0",
  2533 => x"fbdfc287",
  2534 => x"f478c048",
  2535 => x"87e8f28e",
  2536 => x"5c5b5e0e",
  2537 => x"711e0e5d",
  2538 => x"c2cbc44c",
  2539 => x"cdc149bf",
  2540 => x"d1c14da1",
  2541 => x"747e6981",
  2542 => x"87cf029c",
  2543 => x"744ba5c4",
  2544 => x"c2cbc47b",
  2545 => x"c7f249bf",
  2546 => x"747b6e87",
  2547 => x"87c4059c",
  2548 => x"87c24bc0",
  2549 => x"49734bc1",
  2550 => x"d487c8f2",
  2551 => x"87c90266",
  2552 => x"e4cbc149",
  2553 => x"c24a7087",
  2554 => x"c24ac087",
  2555 => x"265affdf",
  2556 => x"0087d5f1",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"1e000000",
  2560 => x"4b711e73",
  2561 => x"4acbc149",
  2562 => x"87c7e9fd",
  2563 => x"721e4a70",
  2564 => x"4afcc049",
  2565 => x"87fbe8fd",
  2566 => x"4a264970",
  2567 => x"714866c8",
  2568 => x"c0497250",
  2569 => x"e8fd4afc",
  2570 => x"4a7187e9",
  2571 => x"c14966c8",
  2572 => x"73517281",
  2573 => x"4acbc149",
  2574 => x"87d7e8fd",
  2575 => x"66c84a71",
  2576 => x"7281c249",
  2577 => x"2687c451",
  2578 => x"264c264d",
  2579 => x"1e4f264b",
  2580 => x"4b711e73",
  2581 => x"c14966c8",
  2582 => x"66cc91cb",
  2583 => x"7349a14a",
  2584 => x"d4c6c14a",
  2585 => x"49a17292",
  2586 => x"7189d6c2",
  2587 => x"87dbff48",
  2588 => x"5c5b5e0e",
  2589 => x"711e0e5d",
  2590 => x"026b974b",
  2591 => x"9787e4c0",
  2592 => x"c0487e6b",
  2593 => x"04a8b7f0",
  2594 => x"486e87d9",
  2595 => x"a8b7f9c0",
  2596 => x"c187d001",
  2597 => x"c0496e83",
  2598 => x"91ca89f0",
  2599 => x"714866d4",
  2600 => x"c087c550",
  2601 => x"87ebc448",
  2602 => x"c0026b97",
  2603 => x"6b9787e9",
  2604 => x"f0c0487e",
  2605 => x"de04a8b7",
  2606 => x"c0486e87",
  2607 => x"01a8b7f9",
  2608 => x"83c187d5",
  2609 => x"f0c0496e",
  2610 => x"9766d489",
  2611 => x"49a14abf",
  2612 => x"714866d4",
  2613 => x"c087c550",
  2614 => x"87f7c348",
  2615 => x"cd026b97",
  2616 => x"496b9787",
  2617 => x"05a9fac0",
  2618 => x"83c187c4",
  2619 => x"48c087c5",
  2620 => x"9787e0c3",
  2621 => x"e7c0026b",
  2622 => x"7e6b9787",
  2623 => x"b7f0c048",
  2624 => x"87dc04a8",
  2625 => x"f9c0486e",
  2626 => x"d301a8b7",
  2627 => x"6e83c187",
  2628 => x"89f0c049",
  2629 => x"66d491ca",
  2630 => x"7184c14c",
  2631 => x"87c57c97",
  2632 => x"eec248c0",
  2633 => x"026b9787",
  2634 => x"9787e4c0",
  2635 => x"c0487e6b",
  2636 => x"04a8b7f0",
  2637 => x"486e87d9",
  2638 => x"a8b7f9c0",
  2639 => x"c187d001",
  2640 => x"c0496e83",
  2641 => x"6c9789f0",
  2642 => x"9749a14a",
  2643 => x"c087c57c",
  2644 => x"87ffc148",
  2645 => x"cd026b97",
  2646 => x"496b9787",
  2647 => x"05a9fac0",
  2648 => x"83c187c4",
  2649 => x"48c087c5",
  2650 => x"9787e8c1",
  2651 => x"e4c0026b",
  2652 => x"4a6b9787",
  2653 => x"aab7f0c0",
  2654 => x"c087da04",
  2655 => x"01aab7f9",
  2656 => x"83c187d3",
  2657 => x"f0c04972",
  2658 => x"d491ca89",
  2659 => x"85c24d66",
  2660 => x"c57d9771",
  2661 => x"c048c087",
  2662 => x"6b9787f9",
  2663 => x"87e4c002",
  2664 => x"487e6b97",
  2665 => x"a8b7f0c0",
  2666 => x"6e87d904",
  2667 => x"b7f9c048",
  2668 => x"87d001a8",
  2669 => x"496e83c1",
  2670 => x"9789f0c0",
  2671 => x"49a14a6d",
  2672 => x"87c47d97",
  2673 => x"87cb48c0",
  2674 => x"c4026b97",
  2675 => x"c248c087",
  2676 => x"2648c187",
  2677 => x"0e87f0f9",
  2678 => x"5d5c5b5e",
  2679 => x"7186f80e",
  2680 => x"4b4cc04d",
  2681 => x"49c2ccc4",
  2682 => x"87ffcbfe",
  2683 => x"b7c04a70",
  2684 => x"f2c204aa",
  2685 => x"02aaca87",
  2686 => x"c087ecc2",
  2687 => x"cf02aae0",
  2688 => x"02aac987",
  2689 => x"aacd87ca",
  2690 => x"ca87c502",
  2691 => x"87c605aa",
  2692 => x"c2029c74",
  2693 => x"e2c087d1",
  2694 => x"87cc05aa",
  2695 => x"b9c14974",
  2696 => x"ffc34c71",
  2697 => x"87fcfe9c",
  2698 => x"c1059c74",
  2699 => x"e1c187e7",
  2700 => x"c804aab7",
  2701 => x"b7fac187",
  2702 => x"d8c106aa",
  2703 => x"b7c1c187",
  2704 => x"87c804aa",
  2705 => x"aab7dac1",
  2706 => x"87c9c106",
  2707 => x"aab7f0c0",
  2708 => x"c087c804",
  2709 => x"06aab7f9",
  2710 => x"c187fac0",
  2711 => x"c002aadb",
  2712 => x"ddc187f3",
  2713 => x"ecc002aa",
  2714 => x"aaedc087",
  2715 => x"87e5c002",
  2716 => x"02aadfc1",
  2717 => x"ecc087df",
  2718 => x"87d902aa",
  2719 => x"02aafdc0",
  2720 => x"fec187d3",
  2721 => x"87cd02aa",
  2722 => x"02aafac0",
  2723 => x"efc087c7",
  2724 => x"cffd05aa",
  2725 => x"b7ffc087",
  2726 => x"c7fd03ab",
  2727 => x"49a37587",
  2728 => x"517283c1",
  2729 => x"7587fdfc",
  2730 => x"51c049a3",
  2731 => x"c403aab7",
  2732 => x"df7ec487",
  2733 => x"059b7387",
  2734 => x"a6c487c7",
  2735 => x"d078c348",
  2736 => x"029c7487",
  2737 => x"7ec187c4",
  2738 => x"7ec087c2",
  2739 => x"6e48a6c4",
  2740 => x"7e66c478",
  2741 => x"8ef8486e",
  2742 => x"0e87ecf5",
  2743 => x"5d5c5b5e",
  2744 => x"c44d710e",
  2745 => x"c04bcacb",
  2746 => x"49f8c04a",
  2747 => x"87e6d7fd",
  2748 => x"ccc41e75",
  2749 => x"fcfd49c2",
  2750 => x"86c487d4",
  2751 => x"c5059870",
  2752 => x"c04cc187",
  2753 => x"49c187ea",
  2754 => x"7087eac0",
  2755 => x"c9059c4c",
  2756 => x"cecbc487",
  2757 => x"87dd49bf",
  2758 => x"9c744c70",
  2759 => x"c487cb05",
  2760 => x"c448cacb",
  2761 => x"78bfdecb",
  2762 => x"cbc487c6",
  2763 => x"78c048ce",
  2764 => x"d2f44874",
  2765 => x"5b5e0e87",
  2766 => x"ff0e5d5c",
  2767 => x"4c7186d4",
  2768 => x"c47e97c0",
  2769 => x"50c048a6",
  2770 => x"c05080c0",
  2771 => x"80c05080",
  2772 => x"80c04d50",
  2773 => x"c080c478",
  2774 => x"c080c478",
  2775 => x"c080c478",
  2776 => x"caccc478",
  2777 => x"87c505bf",
  2778 => x"c3d048c1",
  2779 => x"c2ccc487",
  2780 => x"d078c048",
  2781 => x"f478c080",
  2782 => x"ceccc480",
  2783 => x"c0c378bf",
  2784 => x"78c048e2",
  2785 => x"48decbc4",
  2786 => x"ffc278c0",
  2787 => x"c6f949e2",
  2788 => x"58a6dc87",
  2789 => x"cd02a8c3",
  2790 => x"6e9787d0",
  2791 => x"d8029b4b",
  2792 => x"028bc187",
  2793 => x"8b87f5c1",
  2794 => x"87e4c302",
  2795 => x"c4c7028b",
  2796 => x"c8028b87",
  2797 => x"f1cc87c3",
  2798 => x"48a6c487",
  2799 => x"ffc250c0",
  2800 => x"fec24ae2",
  2801 => x"d2fd49d2",
  2802 => x"987087c5",
  2803 => x"c187c605",
  2804 => x"d5cc7e97",
  2805 => x"e2ffc287",
  2806 => x"d7fec24a",
  2807 => x"eed1fd49",
  2808 => x"05987087",
  2809 => x"97c287c6",
  2810 => x"87fecb7e",
  2811 => x"4ae2ffc2",
  2812 => x"49ddfec2",
  2813 => x"87d7d1fd",
  2814 => x"c0059870",
  2815 => x"97c387c6",
  2816 => x"87e6cb7e",
  2817 => x"4ae2ffc2",
  2818 => x"49e4fec2",
  2819 => x"87ffd0fd",
  2820 => x"cb059870",
  2821 => x"97c487d4",
  2822 => x"87cecb7e",
  2823 => x"486697c4",
  2824 => x"58a6e0c0",
  2825 => x"c1059870",
  2826 => x"a6c887cd",
  2827 => x"c778c048",
  2828 => x"c1056697",
  2829 => x"cbc487cd",
  2830 => x"c002bff6",
  2831 => x"80ff87c7",
  2832 => x"fec050c1",
  2833 => x"e2ffc287",
  2834 => x"eecbc41e",
  2835 => x"fdf6fd49",
  2836 => x"7086c487",
  2837 => x"c8c00298",
  2838 => x"48a6c787",
  2839 => x"c5c050c1",
  2840 => x"48a6c587",
  2841 => x"f9c350c4",
  2842 => x"ccc41efa",
  2843 => x"f9fd49c2",
  2844 => x"86c487f8",
  2845 => x"dc87ccc0",
  2846 => x"a8c14866",
  2847 => x"87c3c005",
  2848 => x"c47e97c0",
  2849 => x"c1486697",
  2850 => x"08a6c480",
  2851 => x"87dac950",
  2852 => x"c048a6d4",
  2853 => x"c47866e0",
  2854 => x"c0486697",
  2855 => x"7058a6e0",
  2856 => x"fbc00598",
  2857 => x"c01eca87",
  2858 => x"e2ffc21e",
  2859 => x"e0d3fd49",
  2860 => x"7086c887",
  2861 => x"a6e0c049",
  2862 => x"0266dc59",
  2863 => x"4887d3c0",
  2864 => x"a8b7e3c1",
  2865 => x"87cac001",
  2866 => x"dc49a5c1",
  2867 => x"c002a966",
  2868 => x"a6c587c8",
  2869 => x"c250c248",
  2870 => x"66dc87ce",
  2871 => x"87c8c24d",
  2872 => x"c14866dc",
  2873 => x"ffc105a8",
  2874 => x"e2ffc287",
  2875 => x"f6fdc24a",
  2876 => x"dacdfd49",
  2877 => x"05987087",
  2878 => x"c087cfc0",
  2879 => x"c048a6e0",
  2880 => x"c478f0e4",
  2881 => x"c178c080",
  2882 => x"ffc287c7",
  2883 => x"fdc24ae2",
  2884 => x"ccfd49fc",
  2885 => x"987087f9",
  2886 => x"87cfc005",
  2887 => x"48a6e0c0",
  2888 => x"78f0e4c0",
  2889 => x"78c180c4",
  2890 => x"c287e6c0",
  2891 => x"c24ae2ff",
  2892 => x"fd49c7fe",
  2893 => x"7087d8cc",
  2894 => x"cfc00598",
  2895 => x"a6e0c087",
  2896 => x"c0e0c048",
  2897 => x"c180c478",
  2898 => x"87c5c078",
  2899 => x"c248a6c5",
  2900 => x"05ac7550",
  2901 => x"c487cec0",
  2902 => x"c048e6cb",
  2903 => x"fc7866e0",
  2904 => x"66e4c080",
  2905 => x"7e97c078",
  2906 => x"486697c4",
  2907 => x"a6c480c1",
  2908 => x"f5c55008",
  2909 => x"a6e8c087",
  2910 => x"e2ffc21e",
  2911 => x"87f0eb49",
  2912 => x"987086c4",
  2913 => x"87c8c005",
  2914 => x"c248a6c5",
  2915 => x"87e3c050",
  2916 => x"6697eac0",
  2917 => x"edc01e49",
  2918 => x"1e496697",
  2919 => x"6697f0c0",
  2920 => x"87ebea49",
  2921 => x"497086c8",
  2922 => x"7181d6c2",
  2923 => x"8066c848",
  2924 => x"c058a6cc",
  2925 => x"f1c47e97",
  2926 => x"6697c487",
  2927 => x"a6e0c048",
  2928 => x"05987058",
  2929 => x"ca87d7c0",
  2930 => x"c21ec01e",
  2931 => x"fd49e2ff",
  2932 => x"c887fece",
  2933 => x"ca497086",
  2934 => x"c45997a6",
  2935 => x"66dc87c2",
  2936 => x"05a8c148",
  2937 => x"c087f9c3",
  2938 => x"c21ea6e8",
  2939 => x"e949e2ff",
  2940 => x"86c487fe",
  2941 => x"c0059870",
  2942 => x"a6c587c8",
  2943 => x"c350c248",
  2944 => x"eac087db",
  2945 => x"1e496697",
  2946 => x"6697edc0",
  2947 => x"f0c01e49",
  2948 => x"e8496697",
  2949 => x"86c887f9",
  2950 => x"97c67e70",
  2951 => x"e0c04866",
  2952 => x"987058a6",
  2953 => x"87e1c005",
  2954 => x"ad49a4c1",
  2955 => x"87edc205",
  2956 => x"bfdecbc4",
  2957 => x"87e5c205",
  2958 => x"d6c2496e",
  2959 => x"c8487181",
  2960 => x"cbc48066",
  2961 => x"d4c258e2",
  2962 => x"4866dc87",
  2963 => x"c205a8c1",
  2964 => x"ad7487cb",
  2965 => x"87cec005",
  2966 => x"d6c2496e",
  2967 => x"c8487181",
  2968 => x"cbc48066",
  2969 => x"b7c158de",
  2970 => x"cec106ad",
  2971 => x"cc486e87",
  2972 => x"e0c08866",
  2973 => x"ad7458a6",
  2974 => x"87cec005",
  2975 => x"66d44970",
  2976 => x"d0487191",
  2977 => x"cbc48066",
  2978 => x"a4c158da",
  2979 => x"c005ad49",
  2980 => x"cbc487d8",
  2981 => x"c005bfde",
  2982 => x"496e87d0",
  2983 => x"c881d6c2",
  2984 => x"48718166",
  2985 => x"cbc488c1",
  2986 => x"66dc58e2",
  2987 => x"9166d449",
  2988 => x"66d04871",
  2989 => x"58a6d480",
  2990 => x"6e87ddc0",
  2991 => x"81d6c249",
  2992 => x"719166d4",
  2993 => x"8066d048",
  2994 => x"c158a6d4",
  2995 => x"c7c005ac",
  2996 => x"d6cbc487",
  2997 => x"7866d048",
  2998 => x"6e48a6cc",
  2999 => x"7e97c078",
  3000 => x"486697c4",
  3001 => x"a6c480c1",
  3002 => x"66d85008",
  3003 => x"02a8c448",
  3004 => x"c587c7c0",
  3005 => x"f2026697",
  3006 => x"97c787d0",
  3007 => x"c8c00566",
  3008 => x"48a6c587",
  3009 => x"f1c050c4",
  3010 => x"05ad7487",
  3011 => x"c487ebc0",
  3012 => x"4abfd6cb",
  3013 => x"bff6cbc4",
  3014 => x"70887248",
  3015 => x"e6cbc44a",
  3016 => x"1e7249bf",
  3017 => x"fd4a0972",
  3018 => x"7087f4cb",
  3019 => x"c44a2649",
  3020 => x"48bfdacb",
  3021 => x"cbc48071",
  3022 => x"b77458e2",
  3023 => x"c5c003ad",
  3024 => x"48a6c587",
  3025 => x"97c550c4",
  3026 => x"c9c00266",
  3027 => x"cecbc487",
  3028 => x"c078c048",
  3029 => x"cbc487c4",
  3030 => x"e8c05dd2",
  3031 => x"cbc41ea6",
  3032 => x"e249bfda",
  3033 => x"86c487d9",
  3034 => x"5ceecbc4",
  3035 => x"486697c5",
  3036 => x"e38ed4ff",
  3037 => x"554187d1",
  3038 => x"004f4944",
  3039 => x"45444f4d",
  3040 => x"33322f31",
  3041 => x"4d003235",
  3042 => x"3145444f",
  3043 => x"3430322f",
  3044 => x"49460038",
  3045 => x"5400454c",
  3046 => x"4b434152",
  3047 => x"45525000",
  3048 => x"00504147",
  3049 => x"45444e49",
  3050 => x"5e0e0058",
  3051 => x"710e5c5b",
  3052 => x"c44cc14b",
  3053 => x"b7bfdacb",
  3054 => x"87d004ab",
  3055 => x"bfdecbc4",
  3056 => x"c701abb7",
  3057 => x"eacbc487",
  3058 => x"87d348bf",
  3059 => x"e4ed4974",
  3060 => x"c484c187",
  3061 => x"b7bfcecb",
  3062 => x"d6ff06ac",
  3063 => x"e148ff87",
  3064 => x"000087e7",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"731e0000",
  3082 => x"4a4b711e",
  3083 => x"ca49721e",
  3084 => x"dec8fd4a",
  3085 => x"26497087",
  3086 => x"7191d04a",
  3087 => x"ca49721e",
  3088 => x"cec8fd4a",
  3089 => x"264a7187",
  3090 => x"49a17249",
  3091 => x"7199ffc3",
  3092 => x"2687c448",
  3093 => x"264c264d",
  3094 => x"1e4f264b",
  3095 => x"4b711e73",
  3096 => x"b7c4494a",
  3097 => x"cf91ca29",
  3098 => x"49a1729a",
  3099 => x"7199ffc3",
  3100 => x"1e87e448",
  3101 => x"4a711e73",
  3102 => x"7087e049",
  3103 => x"059b4b49",
  3104 => x"4bc187c2",
  3105 => x"bfcecbc4",
  3106 => x"c106abb7",
  3107 => x"49734b87",
  3108 => x"7387e2ea",
  3109 => x"87fffe48",
  3110 => x"caf1c41e",
  3111 => x"f1c45997",
  3112 => x"66c448c7",
  3113 => x"5066c850",
  3114 => x"265066cc",
  3115 => x"1e731e4f",
  3116 => x"d0ff4b71",
  3117 => x"78c5c848",
  3118 => x"c148d4ff",
  3119 => x"497378e1",
  3120 => x"2ab7c84a",
  3121 => x"ffc37872",
  3122 => x"ff787199",
  3123 => x"78c448d0",
  3124 => x"1e87c4fe",
  3125 => x"9fc4f2c4",
  3126 => x"d4f1c459",
  3127 => x"2678c148",
  3128 => x"5b5e0e4f",
  3129 => x"4c710e5c",
  3130 => x"c848d0ff",
  3131 => x"d4ff78c5",
  3132 => x"78e4c148",
  3133 => x"4a4966cc",
  3134 => x"729affc3",
  3135 => x"4a66cc78",
  3136 => x"ffc32ac8",
  3137 => x"4b66d09a",
  3138 => x"b27333c7",
  3139 => x"1e717872",
  3140 => x"c5fd4974",
  3141 => x"d0ff87ee",
  3142 => x"2678c448",
  3143 => x"1e87f6fc",
  3144 => x"e0c01e73",
  3145 => x"cbc44bc0",
  3146 => x"c102bfe2",
  3147 => x"f1c487e7",
  3148 => x"c048bfdf",
  3149 => x"c104a8b7",
  3150 => x"cbc487db",
  3151 => x"02abbfe6",
  3152 => x"cbc487d3",
  3153 => x"d049bffe",
  3154 => x"c41e7181",
  3155 => x"fd49eecb",
  3156 => x"c487dde8",
  3157 => x"c41e7386",
  3158 => x"c41ed6cc",
  3159 => x"fd49eecb",
  3160 => x"c887f4e9",
  3161 => x"e6cbc486",
  3162 => x"d602abbf",
  3163 => x"e0c04987",
  3164 => x"cbc489d0",
  3165 => x"7181bffe",
  3166 => x"eecbc41e",
  3167 => x"efe7fd49",
  3168 => x"c886c487",
  3169 => x"731e4966",
  3170 => x"d6ccc41e",
  3171 => x"87d1fd49",
  3172 => x"e1c086c8",
  3173 => x"f0e4c087",
  3174 => x"d6ccc41e",
  3175 => x"eecbc41e",
  3176 => x"f2e8fd49",
  3177 => x"4966d087",
  3178 => x"f0e4c01e",
  3179 => x"d6ccc41e",
  3180 => x"87edfc49",
  3181 => x"defa86d0",
  3182 => x"cbc41e87",
  3183 => x"db05bff6",
  3184 => x"cef1c487",
  3185 => x"c050c148",
  3186 => x"1ecb1e1e",
  3187 => x"c7fb49c2",
  3188 => x"c186cc87",
  3189 => x"87d5fb49",
  3190 => x"87c248c0",
  3191 => x"4f2648c1",
  3192 => x"c41e731e",
  3193 => x"48bfcaf1",
  3194 => x"c006a8c0",
  3195 => x"ebc387e9",
  3196 => x"c049bfc5",
  3197 => x"7087dee3",
  3198 => x"e3c70298",
  3199 => x"c049cd87",
  3200 => x"7087c6e3",
  3201 => x"c9ebc349",
  3202 => x"caf1c459",
  3203 => x"88c148bf",
  3204 => x"58cef1c4",
  3205 => x"c487c9c7",
  3206 => x"bf97cef1",
  3207 => x"05aac24a",
  3208 => x"c487cac3",
  3209 => x"48bfdbf1",
  3210 => x"bfcecbc4",
  3211 => x"c906a8b7",
  3212 => x"cef1c487",
  3213 => x"c650c048",
  3214 => x"f1c487e6",
  3215 => x"02bf97d9",
  3216 => x"c487ddc6",
  3217 => x"05bff6cb",
  3218 => x"f1c487da",
  3219 => x"50c148ce",
  3220 => x"cb1e1ec0",
  3221 => x"f849c21e",
  3222 => x"86cc87fe",
  3223 => x"f2f949c1",
  3224 => x"87fcc587",
  3225 => x"48d9f1c4",
  3226 => x"cbc450c0",
  3227 => x"cd02bfe2",
  3228 => x"c01ec187",
  3229 => x"fa49c0e0",
  3230 => x"86c487e5",
  3231 => x"f1c487d5",
  3232 => x"c448bfdf",
  3233 => x"b7bfdacb",
  3234 => x"c6c004a8",
  3235 => x"cff1c487",
  3236 => x"c450c048",
  3237 => x"48bfe3f1",
  3238 => x"f1c488c1",
  3239 => x"987058e7",
  3240 => x"87cbc005",
  3241 => x"eaf849c0",
  3242 => x"cef1c487",
  3243 => x"c450c048",
  3244 => x"48bfdff1",
  3245 => x"f1c480c1",
  3246 => x"cbc458e3",
  3247 => x"a8b7bfde",
  3248 => x"87dcc404",
  3249 => x"bfdbf1c4",
  3250 => x"c480c148",
  3251 => x"7058dff1",
  3252 => x"87e1e149",
  3253 => x"48cff1c4",
  3254 => x"cbc450c1",
  3255 => x"1e49bfd6",
  3256 => x"49eecbc4",
  3257 => x"87c8e2fd",
  3258 => x"f3c386c4",
  3259 => x"05aac387",
  3260 => x"c487edc3",
  3261 => x"05bff6cb",
  3262 => x"c487dac0",
  3263 => x"c148cef1",
  3264 => x"1e1ec050",
  3265 => x"49c21ecb",
  3266 => x"cc87cdf6",
  3267 => x"f749c186",
  3268 => x"cbc387c1",
  3269 => x"dff1c487",
  3270 => x"cdf249bf",
  3271 => x"dff1c487",
  3272 => x"daf1c458",
  3273 => x"c105bf97",
  3274 => x"4bc087d5",
  3275 => x"bffbf1c4",
  3276 => x"a8b7c048",
  3277 => x"87c7c104",
  3278 => x"bfe2cbc4",
  3279 => x"87e8c005",
  3280 => x"bfdff1c4",
  3281 => x"dacbc449",
  3282 => x"e4c089bf",
  3283 => x"cbc491f0",
  3284 => x"7181bfd6",
  3285 => x"eecbc41e",
  3286 => x"d3e0fd49",
  3287 => x"c01ec087",
  3288 => x"f649f0e4",
  3289 => x"86c887f9",
  3290 => x"bfdff1c4",
  3291 => x"c480c148",
  3292 => x"c158e3f1",
  3293 => x"fbf1c483",
  3294 => x"06abb7bf",
  3295 => x"c487f9fe",
  3296 => x"c048fbf1",
  3297 => x"dff1c478",
  3298 => x"f1c448bf",
  3299 => x"a8b7bff7",
  3300 => x"87d7c003",
  3301 => x"bfe2cbc4",
  3302 => x"87cfc005",
  3303 => x"bfdbf1c4",
  3304 => x"cecbc448",
  3305 => x"06a8b7bf",
  3306 => x"c487f5c0",
  3307 => x"bf97fff1",
  3308 => x"05a9c149",
  3309 => x"c487d2c0",
  3310 => x"c448dff1",
  3311 => x"78bff3f1",
  3312 => x"48caf1c4",
  3313 => x"c6c078c2",
  3314 => x"cef1c487",
  3315 => x"c450c048",
  3316 => x"bf97fff1",
  3317 => x"05a9c249",
  3318 => x"c087c5c0",
  3319 => x"87f3f349",
  3320 => x"0e87f4f1",
  3321 => x"5d5c5b5e",
  3322 => x"86c4ff0e",
  3323 => x"4ac04b76",
  3324 => x"fc49e0c0",
  3325 => x"ff87dff3",
  3326 => x"c5c848d0",
  3327 => x"48d4ff78",
  3328 => x"c078e2c1",
  3329 => x"c048a6e0",
  3330 => x"48d4ff78",
  3331 => x"e4c078c0",
  3332 => x"e0c049a6",
  3333 => x"51688166",
  3334 => x"4866e0c0",
  3335 => x"e4c080c1",
  3336 => x"b7cc58a6",
  3337 => x"e0ff04a8",
  3338 => x"48d0ff87",
  3339 => x"e4c078c4",
  3340 => x"9c4c6697",
  3341 => x"87f3c002",
  3342 => x"c0028cc3",
  3343 => x"8cc587fe",
  3344 => x"87e5c602",
  3345 => x"c8028ccd",
  3346 => x"c3c387e9",
  3347 => x"fbc8028c",
  3348 => x"028cc187",
  3349 => x"8c87d2cc",
  3350 => x"87c9d002",
  3351 => x"d0028cc3",
  3352 => x"8cc187da",
  3353 => x"87f8c102",
  3354 => x"f587ccd4",
  3355 => x"987087cb",
  3356 => x"87ddd402",
  3357 => x"f4f049c0",
  3358 => x"87d5d487",
  3359 => x"c17e97d2",
  3360 => x"c0c248a6",
  3361 => x"50f0c150",
  3362 => x"f1c480c1",
  3363 => x"50bf97c6",
  3364 => x"50ca80c4",
  3365 => x"f1c480c4",
  3366 => x"50bf97c7",
  3367 => x"97c8f1c4",
  3368 => x"f1c450bf",
  3369 => x"50bf97c9",
  3370 => x"48c9f1c4",
  3371 => x"f1c450c0",
  3372 => x"f1c448c8",
  3373 => x"50bf97c9",
  3374 => x"48c7f1c4",
  3375 => x"97c8f1c4",
  3376 => x"f1c450bf",
  3377 => x"f1c448c6",
  3378 => x"50bf97c7",
  3379 => x"1ed21ec1",
  3380 => x"f049a6ca",
  3381 => x"86c887cb",
  3382 => x"d0ef49c0",
  3383 => x"87f1d287",
  3384 => x"7087d6f3",
  3385 => x"e8d20298",
  3386 => x"97e5c087",
  3387 => x"e4c04866",
  3388 => x"987058a6",
  3389 => x"4887da02",
  3390 => x"e4c088c1",
  3391 => x"987058a6",
  3392 => x"87edc002",
  3393 => x"c088c148",
  3394 => x"7058a6e4",
  3395 => x"ebc10298",
  3396 => x"7e97c287",
  3397 => x"c248a6c1",
  3398 => x"50c150c0",
  3399 => x"bfcecbc4",
  3400 => x"87c2ec49",
  3401 => x"5008a6c3",
  3402 => x"48a6e0c0",
  3403 => x"e2c278c2",
  3404 => x"cacbc487",
  3405 => x"d6c249bf",
  3406 => x"a6f0c081",
  3407 => x"caff711e",
  3408 => x"86c487fd",
  3409 => x"a6c17e97",
  3410 => x"50c0c248",
  3411 => x"6697f0c0",
  3412 => x"87d2eb49",
  3413 => x"5008a6c2",
  3414 => x"6697f1c0",
  3415 => x"87c6eb49",
  3416 => x"5008a6c3",
  3417 => x"6697f2c0",
  3418 => x"87faea49",
  3419 => x"5008a6c4",
  3420 => x"c048a6c5",
  3421 => x"c480da50",
  3422 => x"87d7c178",
  3423 => x"6697e6c0",
  3424 => x"87efeb49",
  3425 => x"bfdacbc4",
  3426 => x"81d6c249",
  3427 => x"1ea6f0c0",
  3428 => x"eac9ff71",
  3429 => x"9786c487",
  3430 => x"48a6c17e",
  3431 => x"c050c0c2",
  3432 => x"496697f0",
  3433 => x"c287ffe9",
  3434 => x"c05008a6",
  3435 => x"496697f1",
  3436 => x"c387f3e9",
  3437 => x"c05008a6",
  3438 => x"496697f2",
  3439 => x"c487e7e9",
  3440 => x"c45008a6",
  3441 => x"49bfe2cb",
  3442 => x"a6c931c2",
  3443 => x"db485997",
  3444 => x"c178c480",
  3445 => x"66e4c01e",
  3446 => x"49a6ca1e",
  3447 => x"c887c2ec",
  3448 => x"eb49c086",
  3449 => x"e8ce87c7",
  3450 => x"87cdef87",
  3451 => x"ce029870",
  3452 => x"e5c087df",
  3453 => x"d0496697",
  3454 => x"97e6c031",
  3455 => x"32c84a66",
  3456 => x"e7c0b172",
  3457 => x"b14a6697",
  3458 => x"ffc74d71",
  3459 => x"c09dffff",
  3460 => x"026697e8",
  3461 => x"4887c8c0",
  3462 => x"58a6e4c0",
  3463 => x"c087c7c0",
  3464 => x"c448a6e0",
  3465 => x"497578c0",
  3466 => x"c487ffe5",
  3467 => x"c458dff1",
  3468 => x"c048caf1",
  3469 => x"e3f1c478",
  3470 => x"e3f1c45d",
  3471 => x"66e0c048",
  3472 => x"c4497578",
  3473 => x"89bfdacb",
  3474 => x"bfe6cbc4",
  3475 => x"d6cbc491",
  3476 => x"1e7181bf",
  3477 => x"49eecbc4",
  3478 => x"87d4d4fd",
  3479 => x"f1c486c4",
  3480 => x"78c048ef",
  3481 => x"48d9f1c4",
  3482 => x"f1c450c1",
  3483 => x"50c248ce",
  3484 => x"c087decc",
  3485 => x"026697e8",
  3486 => x"c487c9c0",
  3487 => x"c148d8f1",
  3488 => x"87cdcc50",
  3489 => x"e4e849c0",
  3490 => x"87c5cc87",
  3491 => x"7087eaec",
  3492 => x"fccb0298",
  3493 => x"97edc087",
  3494 => x"c3484966",
  3495 => x"e4c098c0",
  3496 => x"987058a6",
  3497 => x"87dcc002",
  3498 => x"88c0c148",
  3499 => x"58a6e4c0",
  3500 => x"c0029870",
  3501 => x"c14887e9",
  3502 => x"e4c088c0",
  3503 => x"987058a6",
  3504 => x"87c7c102",
  3505 => x"6697e7c0",
  3506 => x"c031d049",
  3507 => x"4a6697e8",
  3508 => x"b17232c8",
  3509 => x"6697e9c0",
  3510 => x"b5714d4a",
  3511 => x"c087f9c0",
  3512 => x"496697e8",
  3513 => x"7087f4e5",
  3514 => x"ebc01e49",
  3515 => x"e5496697",
  3516 => x"497087e9",
  3517 => x"97eec01e",
  3518 => x"dee54966",
  3519 => x"494a7087",
  3520 => x"87cbc5ff",
  3521 => x"4d7086c8",
  3522 => x"c087cdc0",
  3523 => x"496697e6",
  3524 => x"c487e0e5",
  3525 => x"4dbfdacb",
  3526 => x"48caf1c4",
  3527 => x"f1c478c0",
  3528 => x"49755de3",
  3529 => x"c487c3e2",
  3530 => x"c458dff1",
  3531 => x"c45df7f1",
  3532 => x"c448f7f1",
  3533 => x"78bfcacb",
  3534 => x"48fff1c4",
  3535 => x"6697e5c0",
  3536 => x"fbf1c450",
  3537 => x"c478c148",
  3538 => x"bf97fff1",
  3539 => x"c0059949",
  3540 => x"f1c487c9",
  3541 => x"50c448ce",
  3542 => x"c487c6c0",
  3543 => x"c348cef1",
  3544 => x"e549c050",
  3545 => x"e8c887ed",
  3546 => x"87cde987",
  3547 => x"c8029870",
  3548 => x"edc087df",
  3549 => x"48496697",
  3550 => x"c098c0c3",
  3551 => x"7058a6e4",
  3552 => x"dcc00298",
  3553 => x"c0c14887",
  3554 => x"a6e4c088",
  3555 => x"02987058",
  3556 => x"4887e9c0",
  3557 => x"c088c0c1",
  3558 => x"7058a6e4",
  3559 => x"c7c10298",
  3560 => x"97e7c087",
  3561 => x"31d04966",
  3562 => x"6697e8c0",
  3563 => x"7232c84a",
  3564 => x"97e9c0b1",
  3565 => x"714d4a66",
  3566 => x"87eec1b5",
  3567 => x"6697e8c0",
  3568 => x"87d7e249",
  3569 => x"c01e4970",
  3570 => x"496697eb",
  3571 => x"7087cce2",
  3572 => x"eec01e49",
  3573 => x"e2496697",
  3574 => x"4a7087c1",
  3575 => x"eec1ff49",
  3576 => x"7086c887",
  3577 => x"87c2c14d",
  3578 => x"6697e6c0",
  3579 => x"87ebe149",
  3580 => x"c0484970",
  3581 => x"7058a6e4",
  3582 => x"c6c00598",
  3583 => x"a6e0c087",
  3584 => x"c078c148",
  3585 => x"c44866e0",
  3586 => x"b7bfcecb",
  3587 => x"ccc006a8",
  3588 => x"a6e0c087",
  3589 => x"cacbc448",
  3590 => x"c9c078bf",
  3591 => x"a6e0c087",
  3592 => x"decbc448",
  3593 => x"e0c078bf",
  3594 => x"f1c44d66",
  3595 => x"e5c048ff",
  3596 => x"c4506697",
  3597 => x"c45dfbf1",
  3598 => x"bf97fff1",
  3599 => x"c0059949",
  3600 => x"f1c487c9",
  3601 => x"50c048ce",
  3602 => x"c487c6c0",
  3603 => x"c348cef1",
  3604 => x"fff1c450",
  3605 => x"c249bf97",
  3606 => x"f4c402a9",
  3607 => x"e149c087",
  3608 => x"ecc487cb",
  3609 => x"87d1e587",
  3610 => x"c4029870",
  3611 => x"f1c487e3",
  3612 => x"50c448ce",
  3613 => x"f4e049c0",
  3614 => x"87d5c487",
  3615 => x"7087fae4",
  3616 => x"ccc40298",
  3617 => x"dff1c487",
  3618 => x"cbc448bf",
  3619 => x"c088bfda",
  3620 => x"ca58a6e4",
  3621 => x"a6c17e97",
  3622 => x"50c0c248",
  3623 => x"97cef1c4",
  3624 => x"f7c048bf",
  3625 => x"a8c458a6",
  3626 => x"87c9c005",
  3627 => x"48a6f3c0",
  3628 => x"e1c078c2",
  3629 => x"66f3c087",
  3630 => x"05a8c348",
  3631 => x"c087c9c0",
  3632 => x"c048a6f7",
  3633 => x"87c6c078",
  3634 => x"48a6f7c0",
  3635 => x"f3c078c3",
  3636 => x"f7c048a6",
  3637 => x"a6c27866",
  3638 => x"66f3c048",
  3639 => x"c450c050",
  3640 => x"49bfdbf1",
  3641 => x"dcff81c1",
  3642 => x"a6c487fc",
  3643 => x"f1c45008",
  3644 => x"ff49bfdb",
  3645 => x"c587efdc",
  3646 => x"c05008a6",
  3647 => x"1e4ba6f0",
  3648 => x"4966e4c0",
  3649 => x"87f7fbfe",
  3650 => x"6697f4c0",
  3651 => x"d5dcff49",
  3652 => x"08a6ca87",
  3653 => x"97f5c050",
  3654 => x"dcff4966",
  3655 => x"a6cb87c8",
  3656 => x"f6c05008",
  3657 => x"ff496697",
  3658 => x"cc87fbdb",
  3659 => x"735008a6",
  3660 => x"dff1c41e",
  3661 => x"fbfe49bf",
  3662 => x"f8c087c5",
  3663 => x"ff496697",
  3664 => x"d187e3db",
  3665 => x"c05008a6",
  3666 => x"496697f9",
  3667 => x"87d6dbff",
  3668 => x"5008a6d2",
  3669 => x"6697fac0",
  3670 => x"c9dbff49",
  3671 => x"08a6d387",
  3672 => x"ca1ec150",
  3673 => x"49a6d21e",
  3674 => x"87f5ddff",
  3675 => x"49c086d0",
  3676 => x"87f9dcff",
  3677 => x"c087dac0",
  3678 => x"e0c01e1e",
  3679 => x"ff49c51e",
  3680 => x"cc87d5dc",
  3681 => x"d4f1c486",
  3682 => x"c178c048",
  3683 => x"dcdcff49",
  3684 => x"8ec4ff87",
  3685 => x"87fbdaff",
  3686 => x"ff86f41e",
  3687 => x"c5c848d0",
  3688 => x"48d4ff78",
  3689 => x"c078e3c1",
  3690 => x"48d4ff4a",
  3691 => x"497678c0",
  3692 => x"51688172",
  3693 => x"b7ca82c1",
  3694 => x"87ed04aa",
  3695 => x"c448d0ff",
  3696 => x"268ef478",
  3697 => x"f1c41e4f",
  3698 => x"50c148d9",
  3699 => x"c41e4f26",
  3700 => x"c048caf1",
  3701 => x"dbf1c478",
  3702 => x"7840c048",
  3703 => x"48e7f1c4",
  3704 => x"f1c478c0",
  3705 => x"50c148cf",
  3706 => x"bff6cbc4",
  3707 => x"c087c402",
  3708 => x"c187c249",
  3709 => x"d2f1c449",
  3710 => x"f1c45997",
  3711 => x"40c048eb",
  3712 => x"d4f1c478",
  3713 => x"5040c048",
  3714 => x"f3f1c450",
  3715 => x"7840c048",
  3716 => x"48fff1c4",
  3717 => x"789f50c0",
  3718 => x"48daf1c4",
  3719 => x"4f2650c1",
  3720 => x"ff1e731e",
  3721 => x"c5c848d0",
  3722 => x"48d4ff78",
  3723 => x"6878e0c1",
  3724 => x"99ffc349",
  3725 => x"c448d0ff",
  3726 => x"494b7178",
  3727 => x"c30299c1",
  3728 => x"87dfe687",
  3729 => x"99c24973",
  3730 => x"fd87c302",
  3731 => x"497387ca",
  3732 => x"c30299c4",
  3733 => x"87edfd87",
  3734 => x"99c84973",
  3735 => x"fd87d602",
  3736 => x"d0ff87ec",
  3737 => x"78c5c848",
  3738 => x"c148d4ff",
  3739 => x"78c078e6",
  3740 => x"c448d0ff",
  3741 => x"d0497378",
  3742 => x"def1c499",
  3743 => x"ddff5997",
  3744 => x"f1c487de",
  3745 => x"d702bfd4",
  3746 => x"caf1c487",
  3747 => x"87d005bf",
  3748 => x"9fc0f2c4",
  3749 => x"d8ff49bf",
  3750 => x"f1c487d3",
  3751 => x"78c048d4",
  3752 => x"97d8f1c4",
  3753 => x"87d902bf",
  3754 => x"c848d0ff",
  3755 => x"d4ff78c5",
  3756 => x"78e5c148",
  3757 => x"d0ff78c0",
  3758 => x"c478c448",
  3759 => x"c048d8f1",
  3760 => x"d2d6ff50",
  3761 => x"00000087",
  3762 => x"4a711e00",
  3763 => x"49bfc8ff",
  3764 => x"2648a172",
  3765 => x"c8ff1e4f",
  3766 => x"c0fe89bf",
  3767 => x"c0c0c0c0",
  3768 => x"87c401a9",
  3769 => x"87c24ac0",
  3770 => x"48724ac1",
  3771 => x"5e0e4f26",
  3772 => x"0e5d5c5b",
  3773 => x"d4ff4b71",
  3774 => x"4866d04c",
  3775 => x"49d678c0",
  3776 => x"87dfcffe",
  3777 => x"6c7cffc3",
  3778 => x"99ffc349",
  3779 => x"c3494d71",
  3780 => x"e0c199f0",
  3781 => x"87cb05a9",
  3782 => x"6c7cffc3",
  3783 => x"d098c348",
  3784 => x"c3780866",
  3785 => x"4a6c7cff",
  3786 => x"c331c849",
  3787 => x"4a6c7cff",
  3788 => x"4972b271",
  3789 => x"ffc331c8",
  3790 => x"714a6c7c",
  3791 => x"c84972b2",
  3792 => x"7cffc331",
  3793 => x"b2714a6c",
  3794 => x"c048d0ff",
  3795 => x"9b7378e0",
  3796 => x"7287c202",
  3797 => x"2648757b",
  3798 => x"264c264d",
  3799 => x"1e4f264b",
  3800 => x"5e0e4f26",
  3801 => x"f80e5c5b",
  3802 => x"c81e7686",
  3803 => x"fdfd49a6",
  3804 => x"7086c487",
  3805 => x"c0486e4b",
  3806 => x"f0c201a8",
  3807 => x"c34a7387",
  3808 => x"d0c19af0",
  3809 => x"87c702aa",
  3810 => x"05aae0c1",
  3811 => x"7387dec2",
  3812 => x"0299c849",
  3813 => x"c6ff87c3",
  3814 => x"c34c7387",
  3815 => x"05acc29c",
  3816 => x"c487c2c1",
  3817 => x"31c94966",
  3818 => x"66c41e71",
  3819 => x"c492d44a",
  3820 => x"7249c2f2",
  3821 => x"f7fefc81",
  3822 => x"fe49d887",
  3823 => x"c887e4cc",
  3824 => x"f9c31ec0",
  3825 => x"dbfc49fa",
  3826 => x"d0ff87d0",
  3827 => x"78e0c048",
  3828 => x"1efaf9c3",
  3829 => x"d44a66cc",
  3830 => x"c2f2c492",
  3831 => x"fc817249",
  3832 => x"cc87cafd",
  3833 => x"05acc186",
  3834 => x"c487c2c1",
  3835 => x"31c94966",
  3836 => x"66c41e71",
  3837 => x"c492d44a",
  3838 => x"7249c2f2",
  3839 => x"effdfc81",
  3840 => x"faf9c387",
  3841 => x"4a66c81e",
  3842 => x"f2c492d4",
  3843 => x"817249c2",
  3844 => x"87d6fbfc",
  3845 => x"cbfe49d7",
  3846 => x"c0c887c9",
  3847 => x"faf9c31e",
  3848 => x"dfd9fc49",
  3849 => x"ff86cc87",
  3850 => x"e0c048d0",
  3851 => x"fc8ef878",
  3852 => x"5e0e87e7",
  3853 => x"0e5d5c5b",
  3854 => x"ff4d711e",
  3855 => x"66d44cd4",
  3856 => x"b7c3487e",
  3857 => x"87c506a8",
  3858 => x"e2c148c0",
  3859 => x"fd497587",
  3860 => x"7587dbd1",
  3861 => x"4b66c41e",
  3862 => x"f2c493d4",
  3863 => x"497383c2",
  3864 => x"87eaf6fc",
  3865 => x"4b6b83c8",
  3866 => x"c848d0ff",
  3867 => x"7cdd78e1",
  3868 => x"ffc34973",
  3869 => x"737c7199",
  3870 => x"29b7c849",
  3871 => x"7199ffc3",
  3872 => x"d049737c",
  3873 => x"ffc329b7",
  3874 => x"737c7199",
  3875 => x"29b7d849",
  3876 => x"7cc07c71",
  3877 => x"7c7c7c7c",
  3878 => x"7c7c7c7c",
  3879 => x"c07c7c7c",
  3880 => x"66c478e0",
  3881 => x"fe49dc1e",
  3882 => x"c887ddc9",
  3883 => x"26487386",
  3884 => x"0e87e4fa",
  3885 => x"5d5c5b5e",
  3886 => x"7e711e0e",
  3887 => x"6e4bd4ff",
  3888 => x"d6f2c41e",
  3889 => x"c5f5fc49",
  3890 => x"7086c487",
  3891 => x"c3029d4d",
  3892 => x"f2c487c3",
  3893 => x"6e4cbfde",
  3894 => x"d1cffd49",
  3895 => x"48d0ff87",
  3896 => x"c178c5c8",
  3897 => x"4ac07bd6",
  3898 => x"82c17b15",
  3899 => x"aab7e0c0",
  3900 => x"ff87f504",
  3901 => x"78c448d0",
  3902 => x"c178c5c8",
  3903 => x"7bc17bd3",
  3904 => x"9c7478c4",
  3905 => x"87fcc102",
  3906 => x"7efaf9c3",
  3907 => x"8c4dc0c8",
  3908 => x"03acb7c0",
  3909 => x"c0c887c6",
  3910 => x"4cc04da4",
  3911 => x"97ebc6c4",
  3912 => x"99d049bf",
  3913 => x"c087d202",
  3914 => x"d6f2c41e",
  3915 => x"f9f6fc49",
  3916 => x"7086c487",
  3917 => x"efc04a49",
  3918 => x"faf9c387",
  3919 => x"d6f2c41e",
  3920 => x"e5f6fc49",
  3921 => x"7086c487",
  3922 => x"d0ff4a49",
  3923 => x"78c5c848",
  3924 => x"6e7bd4c1",
  3925 => x"6e7bbf97",
  3926 => x"7080c148",
  3927 => x"058dc17e",
  3928 => x"ff87f0ff",
  3929 => x"78c448d0",
  3930 => x"c5059a72",
  3931 => x"c048c087",
  3932 => x"1ec187e5",
  3933 => x"49d6f2c4",
  3934 => x"87cdf4fc",
  3935 => x"9c7486c4",
  3936 => x"87c4fe05",
  3937 => x"c848d0ff",
  3938 => x"d3c178c5",
  3939 => x"c47bc07b",
  3940 => x"c248c178",
  3941 => x"2648c087",
  3942 => x"4c264d26",
  3943 => x"4f264b26",
  3944 => x"5c5b5e0e",
  3945 => x"cc4b710e",
  3946 => x"87dd0266",
  3947 => x"8cf0c04c",
  3948 => x"7487dd02",
  3949 => x"028ac14a",
  3950 => x"028a87d6",
  3951 => x"028a87d2",
  3952 => x"8ad087ce",
  3953 => x"df87db02",
  3954 => x"fb497387",
  3955 => x"87d887e5",
  3956 => x"49c01e74",
  3957 => x"7487dbf9",
  3958 => x"f949731e",
  3959 => x"86c887d4",
  3960 => x"497387c6",
  3961 => x"87ddd0fd",
  3962 => x"0087effe",
  3963 => x"faf8c31e",
  3964 => x"b9c149bf",
  3965 => x"59fef8c3",
  3966 => x"c348d4ff",
  3967 => x"d0ff78ff",
  3968 => x"78e1c848",
  3969 => x"c148d4ff",
  3970 => x"7131c478",
  3971 => x"48d0ff78",
  3972 => x"2678e0c0",
  3973 => x"f8c31e4f",
  3974 => x"f2c41eee",
  3975 => x"effc49d6",
  3976 => x"86c487ec",
  3977 => x"c3029870",
  3978 => x"87c0ff87",
  3979 => x"35314f26",
  3980 => x"205a484b",
  3981 => x"46432020",
  3982 => x"00000047",
  3983 => x"9f1a0000",
  3984 => x"14111258",
  3985 => x"231c1b1d",
  3986 => x"595aa74a",
  3987 => x"f2f59491",
  3988 => x"f2f5f4eb",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
