//`define DEMISTIFY_NO_MEMCARD
//`define DEMISTIFY_NO_YPBPR
//`define VRAM32 1
//`define CLK_SPEED 96000
`define DEMISTIFY
`define VIVADO
`define NO_CD
`define I2S_AUDIO 1
`define VGA_8BIT 1
