
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"ec",x"f2",x"c4",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"ec",x"f2",x"c4"),
    14 => (x"48",x"d4",x"f9",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e3",x"eb"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"48",x"12",x"1e",x"72"),
    21 => (x"87",x"c4",x"02",x"11"),
    22 => (x"87",x"f6",x"02",x"88"),
    23 => (x"4f",x"26",x"4a",x"26"),
    24 => (x"73",x"1e",x"72",x"1e"),
    25 => (x"11",x"48",x"12",x"1e"),
    26 => (x"4b",x"87",x"ca",x"02"),
    27 => (x"9b",x"98",x"df",x"c3"),
    28 => (x"f0",x"02",x"88",x"73"),
    29 => (x"26",x"4b",x"26",x"87"),
    30 => (x"1e",x"4f",x"26",x"4a"),
    31 => (x"1e",x"72",x"1e",x"73"),
    32 => (x"ca",x"04",x"8b",x"c1"),
    33 => (x"11",x"48",x"12",x"87"),
    34 => (x"88",x"87",x"c4",x"02"),
    35 => (x"26",x"87",x"f1",x"02"),
    36 => (x"26",x"4b",x"26",x"4a"),
    37 => (x"1e",x"74",x"1e",x"4f"),
    38 => (x"1e",x"72",x"1e",x"73"),
    39 => (x"d0",x"04",x"8b",x"c1"),
    40 => (x"11",x"48",x"12",x"87"),
    41 => (x"4c",x"87",x"ca",x"02"),
    42 => (x"9c",x"98",x"df",x"c3"),
    43 => (x"eb",x"02",x"88",x"74"),
    44 => (x"26",x"4a",x"26",x"87"),
    45 => (x"26",x"4c",x"26",x"4b"),
    46 => (x"48",x"73",x"1e",x"4f"),
    47 => (x"02",x"a9",x"73",x"81"),
    48 => (x"53",x"12",x"87",x"c5"),
    49 => (x"26",x"87",x"f6",x"05"),
    50 => (x"66",x"c4",x"1e",x"4f"),
    51 => (x"12",x"48",x"71",x"4a"),
    52 => (x"87",x"fb",x"05",x"51"),
    53 => (x"73",x"1e",x"4f",x"26"),
    54 => (x"a9",x"73",x"81",x"48"),
    55 => (x"f9",x"53",x"72",x"05"),
    56 => (x"0e",x"4f",x"26",x"87"),
    57 => (x"5d",x"5c",x"5b",x"5e"),
    58 => (x"71",x"86",x"f4",x"0e"),
    59 => (x"48",x"a6",x"c4",x"4d"),
    60 => (x"66",x"dc",x"78",x"c0"),
    61 => (x"48",x"a6",x"c8",x"4b"),
    62 => (x"97",x"15",x"78",x"c0"),
    63 => (x"02",x"6e",x"97",x"7e"),
    64 => (x"13",x"87",x"f0",x"c0"),
    65 => (x"da",x"02",x"9c",x"4c"),
    66 => (x"4a",x"6e",x"97",x"87"),
    67 => (x"aa",x"b7",x"49",x"74"),
    68 => (x"c8",x"87",x"c9",x"05"),
    69 => (x"78",x"c1",x"48",x"a6"),
    70 => (x"87",x"c2",x"4c",x"c0"),
    71 => (x"9c",x"74",x"4c",x"13"),
    72 => (x"c8",x"87",x"e6",x"05"),
    73 => (x"87",x"cb",x"02",x"66"),
    74 => (x"c1",x"48",x"66",x"c4"),
    75 => (x"58",x"a6",x"c8",x"80"),
    76 => (x"c4",x"87",x"ff",x"fe"),
    77 => (x"8e",x"f4",x"48",x"66"),
    78 => (x"4c",x"26",x"4d",x"26"),
    79 => (x"4f",x"26",x"4b",x"26"),
    80 => (x"c1",x"4a",x"71",x"1e"),
    81 => (x"04",x"aa",x"b7",x"c1"),
    82 => (x"c6",x"c1",x"87",x"d9"),
    83 => (x"d2",x"01",x"aa",x"b7"),
    84 => (x"48",x"66",x"c4",x"87"),
    85 => (x"ca",x"05",x"a8",x"d0"),
    86 => (x"c0",x"49",x"72",x"87"),
    87 => (x"48",x"71",x"89",x"f7"),
    88 => (x"c1",x"87",x"ec",x"c0"),
    89 => (x"04",x"aa",x"b7",x"e1"),
    90 => (x"e6",x"c1",x"87",x"d8"),
    91 => (x"d1",x"01",x"aa",x"b7"),
    92 => (x"48",x"66",x"c4",x"87"),
    93 => (x"c9",x"05",x"a8",x"d0"),
    94 => (x"c1",x"49",x"72",x"87"),
    95 => (x"48",x"71",x"89",x"d7"),
    96 => (x"f0",x"c0",x"87",x"cd"),
    97 => (x"aa",x"b7",x"c9",x"8a"),
    98 => (x"ff",x"87",x"c2",x"06"),
    99 => (x"26",x"48",x"72",x"4a"),
   100 => (x"5b",x"5e",x"0e",x"4f"),
   101 => (x"f8",x"0e",x"5d",x"5c"),
   102 => (x"c4",x"7e",x"71",x"86"),
   103 => (x"78",x"c0",x"48",x"a6"),
   104 => (x"a7",x"f9",x"c1",x"4c"),
   105 => (x"49",x"66",x"c4",x"1e"),
   106 => (x"c4",x"87",x"f8",x"fc"),
   107 => (x"6e",x"49",x"70",x"86"),
   108 => (x"97",x"83",x"71",x"4b"),
   109 => (x"ed",x"c0",x"49",x"6b"),
   110 => (x"87",x"c6",x"05",x"a9"),
   111 => (x"c1",x"48",x"a6",x"c4"),
   112 => (x"66",x"d8",x"83",x"78"),
   113 => (x"d8",x"87",x"c5",x"02"),
   114 => (x"0b",x"7b",x"0b",x"66"),
   115 => (x"d3",x"05",x"6b",x"97"),
   116 => (x"02",x"66",x"c4",x"87"),
   117 => (x"4a",x"74",x"87",x"c7"),
   118 => (x"c2",x"8a",x"0a",x"c0"),
   119 => (x"72",x"4a",x"74",x"87"),
   120 => (x"87",x"ef",x"c0",x"48"),
   121 => (x"13",x"1e",x"66",x"dc"),
   122 => (x"87",x"d4",x"fd",x"49"),
   123 => (x"4d",x"70",x"86",x"c4"),
   124 => (x"03",x"ad",x"b7",x"c0"),
   125 => (x"66",x"c4",x"87",x"d4"),
   126 => (x"74",x"87",x"c9",x"02"),
   127 => (x"88",x"08",x"c0",x"48"),
   128 => (x"87",x"c2",x"7e",x"70"),
   129 => (x"48",x"6e",x"7e",x"74"),
   130 => (x"66",x"dc",x"87",x"c9"),
   131 => (x"4c",x"a4",x"75",x"94"),
   132 => (x"f8",x"87",x"ef",x"fe"),
   133 => (x"26",x"4d",x"26",x"8e"),
   134 => (x"26",x"4b",x"26",x"4c"),
   135 => (x"1e",x"00",x"20",x"4f"),
   136 => (x"9a",x"72",x"1e",x"73"),
   137 => (x"87",x"e7",x"c0",x"02"),
   138 => (x"4b",x"c1",x"48",x"c0"),
   139 => (x"d1",x"06",x"a9",x"72"),
   140 => (x"06",x"82",x"72",x"87"),
   141 => (x"83",x"73",x"87",x"c9"),
   142 => (x"f4",x"01",x"a9",x"72"),
   143 => (x"c1",x"87",x"c3",x"87"),
   144 => (x"a9",x"72",x"3a",x"b2"),
   145 => (x"80",x"73",x"89",x"03"),
   146 => (x"2b",x"2a",x"c1",x"07"),
   147 => (x"26",x"87",x"f3",x"05"),
   148 => (x"1e",x"4f",x"26",x"4b"),
   149 => (x"4d",x"c4",x"1e",x"75"),
   150 => (x"04",x"a1",x"b7",x"71"),
   151 => (x"81",x"c1",x"b9",x"ff"),
   152 => (x"72",x"07",x"bd",x"c3"),
   153 => (x"ff",x"04",x"a2",x"b7"),
   154 => (x"c1",x"82",x"c1",x"ba"),
   155 => (x"ee",x"fe",x"07",x"bd"),
   156 => (x"04",x"2d",x"c1",x"87"),
   157 => (x"80",x"c1",x"b8",x"ff"),
   158 => (x"ff",x"04",x"2d",x"07"),
   159 => (x"07",x"81",x"c1",x"b9"),
   160 => (x"4f",x"26",x"4d",x"26"),
   161 => (x"ff",x"48",x"11",x"1e"),
   162 => (x"c4",x"78",x"08",x"d4"),
   163 => (x"88",x"c1",x"48",x"66"),
   164 => (x"70",x"58",x"a6",x"c8"),
   165 => (x"87",x"ed",x"05",x"98"),
   166 => (x"ff",x"1e",x"4f",x"26"),
   167 => (x"ff",x"c3",x"48",x"d4"),
   168 => (x"c4",x"51",x"68",x"78"),
   169 => (x"88",x"c1",x"48",x"66"),
   170 => (x"70",x"58",x"a6",x"c8"),
   171 => (x"87",x"eb",x"05",x"98"),
   172 => (x"73",x"1e",x"4f",x"26"),
   173 => (x"4b",x"d4",x"ff",x"1e"),
   174 => (x"6b",x"7b",x"ff",x"c3"),
   175 => (x"7b",x"ff",x"c3",x"4a"),
   176 => (x"32",x"c8",x"49",x"6b"),
   177 => (x"ff",x"c3",x"b1",x"72"),
   178 => (x"c8",x"4a",x"6b",x"7b"),
   179 => (x"c3",x"b2",x"71",x"31"),
   180 => (x"49",x"6b",x"7b",x"ff"),
   181 => (x"b1",x"72",x"32",x"c8"),
   182 => (x"87",x"c4",x"48",x"71"),
   183 => (x"4c",x"26",x"4d",x"26"),
   184 => (x"4f",x"26",x"4b",x"26"),
   185 => (x"5c",x"5b",x"5e",x"0e"),
   186 => (x"4a",x"71",x"0e",x"5d"),
   187 => (x"72",x"4c",x"d4",x"ff"),
   188 => (x"99",x"ff",x"c3",x"49"),
   189 => (x"f9",x"c3",x"7c",x"71"),
   190 => (x"c8",x"05",x"bf",x"d4"),
   191 => (x"48",x"66",x"d0",x"87"),
   192 => (x"a6",x"d4",x"30",x"c9"),
   193 => (x"49",x"66",x"d0",x"58"),
   194 => (x"ff",x"c3",x"29",x"d8"),
   195 => (x"d0",x"7c",x"71",x"99"),
   196 => (x"29",x"d0",x"49",x"66"),
   197 => (x"71",x"99",x"ff",x"c3"),
   198 => (x"49",x"66",x"d0",x"7c"),
   199 => (x"ff",x"c3",x"29",x"c8"),
   200 => (x"d0",x"7c",x"71",x"99"),
   201 => (x"ff",x"c3",x"49",x"66"),
   202 => (x"72",x"7c",x"71",x"99"),
   203 => (x"c3",x"29",x"d0",x"49"),
   204 => (x"7c",x"71",x"99",x"ff"),
   205 => (x"f0",x"c9",x"4b",x"6c"),
   206 => (x"ff",x"c3",x"4d",x"ff"),
   207 => (x"87",x"d0",x"05",x"ab"),
   208 => (x"6c",x"7c",x"ff",x"c3"),
   209 => (x"02",x"8d",x"c1",x"4b"),
   210 => (x"ff",x"c3",x"87",x"c6"),
   211 => (x"87",x"f0",x"02",x"ab"),
   212 => (x"c7",x"fe",x"48",x"73"),
   213 => (x"49",x"c0",x"1e",x"87"),
   214 => (x"c3",x"48",x"d4",x"ff"),
   215 => (x"81",x"c1",x"78",x"ff"),
   216 => (x"a9",x"b7",x"c8",x"c3"),
   217 => (x"26",x"87",x"f1",x"04"),
   218 => (x"1e",x"73",x"1e",x"4f"),
   219 => (x"f8",x"c4",x"87",x"e7"),
   220 => (x"1e",x"c0",x"4b",x"df"),
   221 => (x"c1",x"f0",x"ff",x"c0"),
   222 => (x"e7",x"fd",x"49",x"f7"),
   223 => (x"c1",x"86",x"c4",x"87"),
   224 => (x"ea",x"c0",x"05",x"a8"),
   225 => (x"48",x"d4",x"ff",x"87"),
   226 => (x"c1",x"78",x"ff",x"c3"),
   227 => (x"c0",x"c0",x"c0",x"c0"),
   228 => (x"e1",x"c0",x"1e",x"c0"),
   229 => (x"49",x"e9",x"c1",x"f0"),
   230 => (x"c4",x"87",x"c9",x"fd"),
   231 => (x"05",x"98",x"70",x"86"),
   232 => (x"d4",x"ff",x"87",x"ca"),
   233 => (x"78",x"ff",x"c3",x"48"),
   234 => (x"87",x"cb",x"48",x"c1"),
   235 => (x"c1",x"87",x"e6",x"fe"),
   236 => (x"fd",x"fe",x"05",x"8b"),
   237 => (x"fc",x"48",x"c0",x"87"),
   238 => (x"73",x"1e",x"87",x"e6"),
   239 => (x"48",x"d4",x"ff",x"1e"),
   240 => (x"d3",x"78",x"ff",x"c3"),
   241 => (x"c0",x"1e",x"c0",x"4b"),
   242 => (x"c1",x"c1",x"f0",x"ff"),
   243 => (x"87",x"d4",x"fc",x"49"),
   244 => (x"98",x"70",x"86",x"c4"),
   245 => (x"ff",x"87",x"ca",x"05"),
   246 => (x"ff",x"c3",x"48",x"d4"),
   247 => (x"cb",x"48",x"c1",x"78"),
   248 => (x"87",x"f1",x"fd",x"87"),
   249 => (x"ff",x"05",x"8b",x"c1"),
   250 => (x"48",x"c0",x"87",x"db"),
   251 => (x"0e",x"87",x"f1",x"fb"),
   252 => (x"0e",x"5c",x"5b",x"5e"),
   253 => (x"fd",x"4c",x"d4",x"ff"),
   254 => (x"ea",x"c6",x"87",x"db"),
   255 => (x"f0",x"e1",x"c0",x"1e"),
   256 => (x"fb",x"49",x"c8",x"c1"),
   257 => (x"86",x"c4",x"87",x"de"),
   258 => (x"c8",x"02",x"a8",x"c1"),
   259 => (x"87",x"ea",x"fe",x"87"),
   260 => (x"e2",x"c1",x"48",x"c0"),
   261 => (x"87",x"da",x"fa",x"87"),
   262 => (x"ff",x"cf",x"49",x"70"),
   263 => (x"ea",x"c6",x"99",x"ff"),
   264 => (x"87",x"c8",x"02",x"a9"),
   265 => (x"c0",x"87",x"d3",x"fe"),
   266 => (x"87",x"cb",x"c1",x"48"),
   267 => (x"c0",x"7c",x"ff",x"c3"),
   268 => (x"f4",x"fc",x"4b",x"f1"),
   269 => (x"02",x"98",x"70",x"87"),
   270 => (x"c0",x"87",x"eb",x"c0"),
   271 => (x"f0",x"ff",x"c0",x"1e"),
   272 => (x"fa",x"49",x"fa",x"c1"),
   273 => (x"86",x"c4",x"87",x"de"),
   274 => (x"d9",x"05",x"98",x"70"),
   275 => (x"7c",x"ff",x"c3",x"87"),
   276 => (x"ff",x"c3",x"49",x"6c"),
   277 => (x"7c",x"7c",x"7c",x"7c"),
   278 => (x"02",x"99",x"c0",x"c1"),
   279 => (x"48",x"c1",x"87",x"c4"),
   280 => (x"48",x"c0",x"87",x"d5"),
   281 => (x"ab",x"c2",x"87",x"d1"),
   282 => (x"c0",x"87",x"c4",x"05"),
   283 => (x"c1",x"87",x"c8",x"48"),
   284 => (x"fd",x"fe",x"05",x"8b"),
   285 => (x"f9",x"48",x"c0",x"87"),
   286 => (x"73",x"1e",x"87",x"e4"),
   287 => (x"d4",x"f9",x"c3",x"1e"),
   288 => (x"c7",x"78",x"c1",x"48"),
   289 => (x"48",x"d0",x"ff",x"4b"),
   290 => (x"c8",x"fb",x"78",x"c2"),
   291 => (x"48",x"d0",x"ff",x"87"),
   292 => (x"1e",x"c0",x"78",x"c3"),
   293 => (x"c1",x"d0",x"e5",x"c0"),
   294 => (x"c7",x"f9",x"49",x"c0"),
   295 => (x"c1",x"86",x"c4",x"87"),
   296 => (x"87",x"c1",x"05",x"a8"),
   297 => (x"05",x"ab",x"c2",x"4b"),
   298 => (x"48",x"c0",x"87",x"c5"),
   299 => (x"c1",x"87",x"f9",x"c0"),
   300 => (x"d0",x"ff",x"05",x"8b"),
   301 => (x"87",x"f7",x"fc",x"87"),
   302 => (x"58",x"d8",x"f9",x"c3"),
   303 => (x"cd",x"05",x"98",x"70"),
   304 => (x"c0",x"1e",x"c1",x"87"),
   305 => (x"d0",x"c1",x"f0",x"ff"),
   306 => (x"87",x"d8",x"f8",x"49"),
   307 => (x"d4",x"ff",x"86",x"c4"),
   308 => (x"78",x"ff",x"c3",x"48"),
   309 => (x"c3",x"87",x"e0",x"c4"),
   310 => (x"ff",x"58",x"dc",x"f9"),
   311 => (x"78",x"c2",x"48",x"d0"),
   312 => (x"c3",x"48",x"d4",x"ff"),
   313 => (x"48",x"c1",x"78",x"ff"),
   314 => (x"0e",x"87",x"f5",x"f7"),
   315 => (x"5d",x"5c",x"5b",x"5e"),
   316 => (x"c3",x"4a",x"71",x"0e"),
   317 => (x"d4",x"ff",x"4d",x"ff"),
   318 => (x"ff",x"7c",x"75",x"4c"),
   319 => (x"c3",x"c4",x"48",x"d0"),
   320 => (x"72",x"7c",x"75",x"78"),
   321 => (x"f0",x"ff",x"c0",x"1e"),
   322 => (x"f7",x"49",x"d8",x"c1"),
   323 => (x"86",x"c4",x"87",x"d6"),
   324 => (x"c5",x"02",x"98",x"70"),
   325 => (x"c0",x"48",x"c0",x"87"),
   326 => (x"7c",x"75",x"87",x"f0"),
   327 => (x"c8",x"7c",x"fe",x"c3"),
   328 => (x"66",x"d4",x"1e",x"c0"),
   329 => (x"87",x"dc",x"f5",x"49"),
   330 => (x"7c",x"75",x"86",x"c4"),
   331 => (x"7c",x"75",x"7c",x"75"),
   332 => (x"4b",x"e0",x"da",x"d8"),
   333 => (x"49",x"6c",x"7c",x"75"),
   334 => (x"87",x"c5",x"05",x"99"),
   335 => (x"f3",x"05",x"8b",x"c1"),
   336 => (x"ff",x"7c",x"75",x"87"),
   337 => (x"78",x"c2",x"48",x"d0"),
   338 => (x"cf",x"f6",x"48",x"c1"),
   339 => (x"d4",x"ff",x"1e",x"87"),
   340 => (x"48",x"d0",x"ff",x"4a"),
   341 => (x"c3",x"78",x"d1",x"c4"),
   342 => (x"89",x"c1",x"7a",x"ff"),
   343 => (x"26",x"87",x"f8",x"05"),
   344 => (x"1e",x"73",x"1e",x"4f"),
   345 => (x"ee",x"c5",x"4b",x"71"),
   346 => (x"ff",x"4a",x"df",x"cd"),
   347 => (x"ff",x"c3",x"48",x"d4"),
   348 => (x"c3",x"48",x"68",x"78"),
   349 => (x"c5",x"02",x"a8",x"fe"),
   350 => (x"05",x"8a",x"c1",x"87"),
   351 => (x"9a",x"72",x"87",x"ed"),
   352 => (x"c0",x"87",x"c5",x"05"),
   353 => (x"87",x"ea",x"c0",x"48"),
   354 => (x"cc",x"02",x"9b",x"73"),
   355 => (x"1e",x"66",x"c8",x"87"),
   356 => (x"c5",x"f4",x"49",x"73"),
   357 => (x"c6",x"86",x"c4",x"87"),
   358 => (x"49",x"66",x"c8",x"87"),
   359 => (x"ff",x"87",x"ee",x"fe"),
   360 => (x"ff",x"c3",x"48",x"d4"),
   361 => (x"9b",x"73",x"78",x"78"),
   362 => (x"ff",x"87",x"c5",x"05"),
   363 => (x"78",x"d0",x"48",x"d0"),
   364 => (x"eb",x"f4",x"48",x"c1"),
   365 => (x"1e",x"73",x"1e",x"87"),
   366 => (x"4b",x"c0",x"4a",x"71"),
   367 => (x"c3",x"48",x"d4",x"ff"),
   368 => (x"d0",x"ff",x"78",x"ff"),
   369 => (x"78",x"c3",x"c4",x"48"),
   370 => (x"c3",x"48",x"d4",x"ff"),
   371 => (x"1e",x"72",x"78",x"ff"),
   372 => (x"c1",x"f0",x"ff",x"c0"),
   373 => (x"cb",x"f4",x"49",x"d1"),
   374 => (x"70",x"86",x"c4",x"87"),
   375 => (x"87",x"cd",x"05",x"98"),
   376 => (x"cc",x"1e",x"c0",x"c8"),
   377 => (x"f8",x"fd",x"49",x"66"),
   378 => (x"70",x"86",x"c4",x"87"),
   379 => (x"48",x"d0",x"ff",x"4b"),
   380 => (x"48",x"73",x"78",x"c2"),
   381 => (x"0e",x"87",x"e9",x"f3"),
   382 => (x"5d",x"5c",x"5b",x"5e"),
   383 => (x"c0",x"1e",x"c0",x"0e"),
   384 => (x"c9",x"c1",x"f0",x"ff"),
   385 => (x"87",x"dc",x"f3",x"49"),
   386 => (x"f9",x"c3",x"1e",x"d2"),
   387 => (x"d0",x"fd",x"49",x"dc"),
   388 => (x"c0",x"86",x"c8",x"87"),
   389 => (x"d2",x"84",x"c1",x"4c"),
   390 => (x"f8",x"04",x"ac",x"b7"),
   391 => (x"dc",x"f9",x"c3",x"87"),
   392 => (x"c3",x"49",x"bf",x"97"),
   393 => (x"c0",x"c1",x"99",x"c0"),
   394 => (x"e7",x"c0",x"05",x"a9"),
   395 => (x"e3",x"f9",x"c3",x"87"),
   396 => (x"d0",x"49",x"bf",x"97"),
   397 => (x"e4",x"f9",x"c3",x"31"),
   398 => (x"c8",x"4a",x"bf",x"97"),
   399 => (x"c3",x"b1",x"72",x"32"),
   400 => (x"bf",x"97",x"e5",x"f9"),
   401 => (x"4c",x"71",x"b1",x"4a"),
   402 => (x"ff",x"ff",x"ff",x"cf"),
   403 => (x"ca",x"84",x"c1",x"9c"),
   404 => (x"87",x"e7",x"c1",x"34"),
   405 => (x"97",x"e5",x"f9",x"c3"),
   406 => (x"31",x"c1",x"49",x"bf"),
   407 => (x"f9",x"c3",x"99",x"c6"),
   408 => (x"4a",x"bf",x"97",x"e6"),
   409 => (x"72",x"2a",x"b7",x"c7"),
   410 => (x"e1",x"f9",x"c3",x"b1"),
   411 => (x"4d",x"4a",x"bf",x"97"),
   412 => (x"f9",x"c3",x"9d",x"cf"),
   413 => (x"4a",x"bf",x"97",x"e2"),
   414 => (x"32",x"ca",x"9a",x"c3"),
   415 => (x"97",x"e3",x"f9",x"c3"),
   416 => (x"33",x"c2",x"4b",x"bf"),
   417 => (x"f9",x"c3",x"b2",x"73"),
   418 => (x"4b",x"bf",x"97",x"e4"),
   419 => (x"c6",x"9b",x"c0",x"c3"),
   420 => (x"b2",x"73",x"2b",x"b7"),
   421 => (x"48",x"c1",x"81",x"c2"),
   422 => (x"49",x"70",x"30",x"71"),
   423 => (x"30",x"75",x"48",x"c1"),
   424 => (x"4c",x"72",x"4d",x"70"),
   425 => (x"94",x"71",x"84",x"c1"),
   426 => (x"ad",x"b7",x"c0",x"c8"),
   427 => (x"c1",x"87",x"cc",x"06"),
   428 => (x"c8",x"2d",x"b7",x"34"),
   429 => (x"01",x"ad",x"b7",x"c0"),
   430 => (x"74",x"87",x"f4",x"ff"),
   431 => (x"87",x"dc",x"f0",x"48"),
   432 => (x"5c",x"5b",x"5e",x"0e"),
   433 => (x"86",x"f8",x"0e",x"5d"),
   434 => (x"48",x"c2",x"c2",x"c4"),
   435 => (x"f9",x"c3",x"78",x"c0"),
   436 => (x"49",x"c0",x"1e",x"fa"),
   437 => (x"c4",x"87",x"de",x"fb"),
   438 => (x"05",x"98",x"70",x"86"),
   439 => (x"48",x"c0",x"87",x"c5"),
   440 => (x"c0",x"87",x"ce",x"c9"),
   441 => (x"c0",x"7e",x"c1",x"4d"),
   442 => (x"49",x"bf",x"f9",x"fe"),
   443 => (x"4a",x"f0",x"fa",x"c3"),
   444 => (x"e6",x"4b",x"c8",x"71"),
   445 => (x"98",x"70",x"87",x"c5"),
   446 => (x"c0",x"87",x"c2",x"05"),
   447 => (x"f5",x"fe",x"c0",x"7e"),
   448 => (x"fb",x"c3",x"49",x"bf"),
   449 => (x"c8",x"71",x"4a",x"cc"),
   450 => (x"87",x"ef",x"e5",x"4b"),
   451 => (x"c2",x"05",x"98",x"70"),
   452 => (x"6e",x"7e",x"c0",x"87"),
   453 => (x"87",x"fd",x"c0",x"02"),
   454 => (x"bf",x"c0",x"c1",x"c4"),
   455 => (x"f8",x"c1",x"c4",x"4d"),
   456 => (x"48",x"7e",x"bf",x"9f"),
   457 => (x"a8",x"ea",x"d6",x"c5"),
   458 => (x"c4",x"87",x"c7",x"05"),
   459 => (x"4d",x"bf",x"c0",x"c1"),
   460 => (x"48",x"6e",x"87",x"ce"),
   461 => (x"a8",x"d5",x"e9",x"ca"),
   462 => (x"c0",x"87",x"c5",x"02"),
   463 => (x"87",x"f1",x"c7",x"48"),
   464 => (x"1e",x"fa",x"f9",x"c3"),
   465 => (x"ec",x"f9",x"49",x"75"),
   466 => (x"70",x"86",x"c4",x"87"),
   467 => (x"87",x"c5",x"05",x"98"),
   468 => (x"dc",x"c7",x"48",x"c0"),
   469 => (x"f5",x"fe",x"c0",x"87"),
   470 => (x"fb",x"c3",x"49",x"bf"),
   471 => (x"c8",x"71",x"4a",x"cc"),
   472 => (x"87",x"d7",x"e4",x"4b"),
   473 => (x"c8",x"05",x"98",x"70"),
   474 => (x"c2",x"c2",x"c4",x"87"),
   475 => (x"da",x"78",x"c1",x"48"),
   476 => (x"f9",x"fe",x"c0",x"87"),
   477 => (x"fa",x"c3",x"49",x"bf"),
   478 => (x"c8",x"71",x"4a",x"f0"),
   479 => (x"87",x"fb",x"e3",x"4b"),
   480 => (x"c0",x"02",x"98",x"70"),
   481 => (x"48",x"c0",x"87",x"c5"),
   482 => (x"c4",x"87",x"e6",x"c6"),
   483 => (x"bf",x"97",x"f8",x"c1"),
   484 => (x"a9",x"d5",x"c1",x"49"),
   485 => (x"87",x"cd",x"c0",x"05"),
   486 => (x"97",x"f9",x"c1",x"c4"),
   487 => (x"ea",x"c2",x"49",x"bf"),
   488 => (x"c5",x"c0",x"02",x"a9"),
   489 => (x"c6",x"48",x"c0",x"87"),
   490 => (x"f9",x"c3",x"87",x"c7"),
   491 => (x"7e",x"bf",x"97",x"fa"),
   492 => (x"a8",x"e9",x"c3",x"48"),
   493 => (x"87",x"ce",x"c0",x"02"),
   494 => (x"eb",x"c3",x"48",x"6e"),
   495 => (x"c5",x"c0",x"02",x"a8"),
   496 => (x"c5",x"48",x"c0",x"87"),
   497 => (x"fa",x"c3",x"87",x"eb"),
   498 => (x"49",x"bf",x"97",x"c5"),
   499 => (x"cc",x"c0",x"05",x"99"),
   500 => (x"c6",x"fa",x"c3",x"87"),
   501 => (x"c2",x"49",x"bf",x"97"),
   502 => (x"c5",x"c0",x"02",x"a9"),
   503 => (x"c5",x"48",x"c0",x"87"),
   504 => (x"fa",x"c3",x"87",x"cf"),
   505 => (x"48",x"bf",x"97",x"c7"),
   506 => (x"58",x"fe",x"c1",x"c4"),
   507 => (x"c1",x"48",x"4c",x"70"),
   508 => (x"c2",x"c2",x"c4",x"88"),
   509 => (x"c8",x"fa",x"c3",x"58"),
   510 => (x"75",x"49",x"bf",x"97"),
   511 => (x"c9",x"fa",x"c3",x"81"),
   512 => (x"c8",x"4a",x"bf",x"97"),
   513 => (x"7e",x"a1",x"72",x"32"),
   514 => (x"48",x"cf",x"c6",x"c4"),
   515 => (x"fa",x"c3",x"78",x"6e"),
   516 => (x"48",x"bf",x"97",x"ca"),
   517 => (x"c4",x"58",x"a6",x"c8"),
   518 => (x"02",x"bf",x"c2",x"c2"),
   519 => (x"c0",x"87",x"d4",x"c2"),
   520 => (x"49",x"bf",x"f5",x"fe"),
   521 => (x"4a",x"cc",x"fb",x"c3"),
   522 => (x"e1",x"4b",x"c8",x"71"),
   523 => (x"98",x"70",x"87",x"cd"),
   524 => (x"87",x"c5",x"c0",x"02"),
   525 => (x"f8",x"c3",x"48",x"c0"),
   526 => (x"fa",x"c1",x"c4",x"87"),
   527 => (x"c6",x"c4",x"4c",x"bf"),
   528 => (x"fa",x"c3",x"5c",x"e3"),
   529 => (x"49",x"bf",x"97",x"df"),
   530 => (x"fa",x"c3",x"31",x"c8"),
   531 => (x"4a",x"bf",x"97",x"de"),
   532 => (x"fa",x"c3",x"49",x"a1"),
   533 => (x"4a",x"bf",x"97",x"e0"),
   534 => (x"a1",x"72",x"32",x"d0"),
   535 => (x"e1",x"fa",x"c3",x"49"),
   536 => (x"d8",x"4a",x"bf",x"97"),
   537 => (x"49",x"a1",x"72",x"32"),
   538 => (x"c4",x"91",x"66",x"c4"),
   539 => (x"81",x"bf",x"cf",x"c6"),
   540 => (x"59",x"d7",x"c6",x"c4"),
   541 => (x"97",x"e7",x"fa",x"c3"),
   542 => (x"32",x"c8",x"4a",x"bf"),
   543 => (x"97",x"e6",x"fa",x"c3"),
   544 => (x"4a",x"a2",x"4b",x"bf"),
   545 => (x"97",x"e8",x"fa",x"c3"),
   546 => (x"33",x"d0",x"4b",x"bf"),
   547 => (x"c3",x"4a",x"a2",x"73"),
   548 => (x"bf",x"97",x"e9",x"fa"),
   549 => (x"d8",x"9b",x"cf",x"4b"),
   550 => (x"4a",x"a2",x"73",x"33"),
   551 => (x"5a",x"db",x"c6",x"c4"),
   552 => (x"bf",x"d7",x"c6",x"c4"),
   553 => (x"74",x"8a",x"c2",x"4a"),
   554 => (x"db",x"c6",x"c4",x"92"),
   555 => (x"78",x"a1",x"72",x"48"),
   556 => (x"c3",x"87",x"ca",x"c1"),
   557 => (x"bf",x"97",x"cc",x"fa"),
   558 => (x"c3",x"31",x"c8",x"49"),
   559 => (x"bf",x"97",x"cb",x"fa"),
   560 => (x"c4",x"49",x"a1",x"4a"),
   561 => (x"c4",x"59",x"ca",x"c2"),
   562 => (x"49",x"bf",x"c6",x"c2"),
   563 => (x"ff",x"c7",x"31",x"c5"),
   564 => (x"c4",x"29",x"c9",x"81"),
   565 => (x"c3",x"59",x"e3",x"c6"),
   566 => (x"bf",x"97",x"d1",x"fa"),
   567 => (x"c3",x"32",x"c8",x"4a"),
   568 => (x"bf",x"97",x"d0",x"fa"),
   569 => (x"c4",x"4a",x"a2",x"4b"),
   570 => (x"82",x"6e",x"92",x"66"),
   571 => (x"5a",x"df",x"c6",x"c4"),
   572 => (x"48",x"d7",x"c6",x"c4"),
   573 => (x"c6",x"c4",x"78",x"c0"),
   574 => (x"a1",x"72",x"48",x"d3"),
   575 => (x"e3",x"c6",x"c4",x"78"),
   576 => (x"d7",x"c6",x"c4",x"48"),
   577 => (x"c6",x"c4",x"78",x"bf"),
   578 => (x"c6",x"c4",x"48",x"e7"),
   579 => (x"c4",x"78",x"bf",x"db"),
   580 => (x"02",x"bf",x"c2",x"c2"),
   581 => (x"74",x"87",x"c9",x"c0"),
   582 => (x"70",x"30",x"c4",x"48"),
   583 => (x"87",x"c9",x"c0",x"7e"),
   584 => (x"bf",x"df",x"c6",x"c4"),
   585 => (x"70",x"30",x"c4",x"48"),
   586 => (x"c6",x"c2",x"c4",x"7e"),
   587 => (x"c1",x"78",x"6e",x"48"),
   588 => (x"26",x"8e",x"f8",x"48"),
   589 => (x"26",x"4c",x"26",x"4d"),
   590 => (x"0e",x"4f",x"26",x"4b"),
   591 => (x"5d",x"5c",x"5b",x"5e"),
   592 => (x"c4",x"4a",x"71",x"0e"),
   593 => (x"02",x"bf",x"c2",x"c2"),
   594 => (x"4b",x"72",x"87",x"cb"),
   595 => (x"4c",x"72",x"2b",x"c7"),
   596 => (x"c9",x"9c",x"ff",x"c1"),
   597 => (x"c8",x"4b",x"72",x"87"),
   598 => (x"c3",x"4c",x"72",x"2b"),
   599 => (x"c6",x"c4",x"9c",x"ff"),
   600 => (x"c0",x"83",x"bf",x"cf"),
   601 => (x"ab",x"bf",x"f1",x"fe"),
   602 => (x"c0",x"87",x"d9",x"02"),
   603 => (x"c3",x"5b",x"f5",x"fe"),
   604 => (x"73",x"1e",x"fa",x"f9"),
   605 => (x"87",x"fd",x"f0",x"49"),
   606 => (x"98",x"70",x"86",x"c4"),
   607 => (x"c0",x"87",x"c5",x"05"),
   608 => (x"87",x"e6",x"c0",x"48"),
   609 => (x"bf",x"c2",x"c2",x"c4"),
   610 => (x"74",x"87",x"d2",x"02"),
   611 => (x"c3",x"91",x"c4",x"49"),
   612 => (x"69",x"81",x"fa",x"f9"),
   613 => (x"ff",x"ff",x"cf",x"4d"),
   614 => (x"cb",x"9d",x"ff",x"ff"),
   615 => (x"c2",x"49",x"74",x"87"),
   616 => (x"fa",x"f9",x"c3",x"91"),
   617 => (x"4d",x"69",x"9f",x"81"),
   618 => (x"c6",x"fe",x"48",x"75"),
   619 => (x"5b",x"5e",x"0e",x"87"),
   620 => (x"1e",x"0e",x"5d",x"5c"),
   621 => (x"1e",x"c0",x"4d",x"71"),
   622 => (x"dc",x"d0",x"49",x"c1"),
   623 => (x"70",x"86",x"c4",x"87"),
   624 => (x"c1",x"02",x"9c",x"4c"),
   625 => (x"c2",x"c4",x"87",x"c2"),
   626 => (x"49",x"75",x"4a",x"ca"),
   627 => (x"87",x"d0",x"da",x"ff"),
   628 => (x"c0",x"02",x"98",x"70"),
   629 => (x"4a",x"74",x"87",x"f2"),
   630 => (x"4b",x"cb",x"49",x"75"),
   631 => (x"87",x"f5",x"da",x"ff"),
   632 => (x"c0",x"02",x"98",x"70"),
   633 => (x"1e",x"c0",x"87",x"e2"),
   634 => (x"c7",x"02",x"9c",x"74"),
   635 => (x"48",x"a6",x"c4",x"87"),
   636 => (x"87",x"c5",x"78",x"c0"),
   637 => (x"c1",x"48",x"a6",x"c4"),
   638 => (x"49",x"66",x"c4",x"78"),
   639 => (x"c4",x"87",x"da",x"cf"),
   640 => (x"9c",x"4c",x"70",x"86"),
   641 => (x"87",x"fe",x"fe",x"05"),
   642 => (x"fc",x"26",x"48",x"74"),
   643 => (x"5e",x"0e",x"87",x"e5"),
   644 => (x"0e",x"5d",x"5c",x"5b"),
   645 => (x"9b",x"4b",x"71",x"1e"),
   646 => (x"c0",x"87",x"c5",x"05"),
   647 => (x"87",x"e5",x"c1",x"48"),
   648 => (x"c0",x"4d",x"a3",x"c8"),
   649 => (x"02",x"66",x"d4",x"7d"),
   650 => (x"66",x"d4",x"87",x"c7"),
   651 => (x"c5",x"05",x"bf",x"97"),
   652 => (x"c1",x"48",x"c0",x"87"),
   653 => (x"66",x"d4",x"87",x"cf"),
   654 => (x"87",x"f1",x"fd",x"49"),
   655 => (x"02",x"9c",x"4c",x"70"),
   656 => (x"dc",x"87",x"c0",x"c1"),
   657 => (x"7d",x"69",x"49",x"a4"),
   658 => (x"c4",x"49",x"a4",x"da"),
   659 => (x"69",x"9f",x"4a",x"a3"),
   660 => (x"c2",x"c2",x"c4",x"7a"),
   661 => (x"87",x"d2",x"02",x"bf"),
   662 => (x"9f",x"49",x"a4",x"d4"),
   663 => (x"ff",x"c0",x"49",x"69"),
   664 => (x"48",x"71",x"99",x"ff"),
   665 => (x"7e",x"70",x"30",x"d0"),
   666 => (x"7e",x"c0",x"87",x"c2"),
   667 => (x"6a",x"48",x"49",x"6e"),
   668 => (x"c0",x"7a",x"70",x"80"),
   669 => (x"49",x"a3",x"cc",x"7b"),
   670 => (x"a3",x"d0",x"79",x"6a"),
   671 => (x"74",x"79",x"c0",x"49"),
   672 => (x"c0",x"87",x"c2",x"48"),
   673 => (x"ea",x"fa",x"26",x"48"),
   674 => (x"5b",x"5e",x"0e",x"87"),
   675 => (x"71",x"0e",x"5d",x"5c"),
   676 => (x"f1",x"fe",x"c0",x"4c"),
   677 => (x"74",x"78",x"ff",x"48"),
   678 => (x"ca",x"c1",x"02",x"9c"),
   679 => (x"49",x"a4",x"c8",x"87"),
   680 => (x"c2",x"c1",x"02",x"69"),
   681 => (x"4a",x"66",x"d0",x"87"),
   682 => (x"d4",x"82",x"49",x"6c"),
   683 => (x"66",x"d0",x"5a",x"a6"),
   684 => (x"c1",x"c4",x"b9",x"4d"),
   685 => (x"ff",x"4a",x"bf",x"fe"),
   686 => (x"71",x"99",x"72",x"ba"),
   687 => (x"e4",x"c0",x"02",x"99"),
   688 => (x"4b",x"a4",x"c4",x"87"),
   689 => (x"f2",x"f9",x"49",x"6b"),
   690 => (x"c4",x"7b",x"70",x"87"),
   691 => (x"49",x"bf",x"fa",x"c1"),
   692 => (x"7c",x"71",x"81",x"6c"),
   693 => (x"c1",x"c4",x"b9",x"75"),
   694 => (x"ff",x"4a",x"bf",x"fe"),
   695 => (x"71",x"99",x"72",x"ba"),
   696 => (x"dc",x"ff",x"05",x"99"),
   697 => (x"f9",x"7c",x"75",x"87"),
   698 => (x"73",x"1e",x"87",x"c9"),
   699 => (x"9b",x"4b",x"71",x"1e"),
   700 => (x"c8",x"87",x"c7",x"02"),
   701 => (x"05",x"69",x"49",x"a3"),
   702 => (x"48",x"c0",x"87",x"c5"),
   703 => (x"c4",x"87",x"eb",x"c0"),
   704 => (x"4a",x"bf",x"d3",x"c6"),
   705 => (x"69",x"49",x"a3",x"c4"),
   706 => (x"c4",x"89",x"c2",x"49"),
   707 => (x"91",x"bf",x"fa",x"c1"),
   708 => (x"c4",x"4a",x"a2",x"71"),
   709 => (x"49",x"bf",x"fe",x"c1"),
   710 => (x"a2",x"71",x"99",x"6b"),
   711 => (x"1e",x"66",x"c8",x"4a"),
   712 => (x"d0",x"ea",x"49",x"72"),
   713 => (x"70",x"86",x"c4",x"87"),
   714 => (x"ca",x"f8",x"48",x"49"),
   715 => (x"1e",x"73",x"1e",x"87"),
   716 => (x"02",x"9b",x"4b",x"71"),
   717 => (x"a3",x"c8",x"87",x"c7"),
   718 => (x"c5",x"05",x"69",x"49"),
   719 => (x"c0",x"48",x"c0",x"87"),
   720 => (x"c6",x"c4",x"87",x"eb"),
   721 => (x"c4",x"4a",x"bf",x"d3"),
   722 => (x"49",x"69",x"49",x"a3"),
   723 => (x"c1",x"c4",x"89",x"c2"),
   724 => (x"71",x"91",x"bf",x"fa"),
   725 => (x"c1",x"c4",x"4a",x"a2"),
   726 => (x"6b",x"49",x"bf",x"fe"),
   727 => (x"4a",x"a2",x"71",x"99"),
   728 => (x"72",x"1e",x"66",x"c8"),
   729 => (x"87",x"c3",x"e6",x"49"),
   730 => (x"49",x"70",x"86",x"c4"),
   731 => (x"87",x"c7",x"f7",x"48"),
   732 => (x"5c",x"5b",x"5e",x"0e"),
   733 => (x"71",x"1e",x"0e",x"5d"),
   734 => (x"4c",x"66",x"d4",x"4b"),
   735 => (x"9b",x"73",x"2c",x"c9"),
   736 => (x"87",x"cf",x"c1",x"02"),
   737 => (x"69",x"49",x"a3",x"c8"),
   738 => (x"87",x"c7",x"c1",x"02"),
   739 => (x"d4",x"4d",x"a3",x"d0"),
   740 => (x"c1",x"c4",x"7d",x"66"),
   741 => (x"ff",x"49",x"bf",x"fe"),
   742 => (x"99",x"4a",x"6b",x"b9"),
   743 => (x"03",x"ac",x"71",x"7e"),
   744 => (x"7b",x"c0",x"87",x"cd"),
   745 => (x"4a",x"a3",x"cc",x"7d"),
   746 => (x"6a",x"49",x"a3",x"c4"),
   747 => (x"72",x"87",x"c2",x"79"),
   748 => (x"02",x"9c",x"74",x"8c"),
   749 => (x"1e",x"49",x"87",x"dd"),
   750 => (x"cc",x"fb",x"49",x"73"),
   751 => (x"d4",x"86",x"c4",x"87"),
   752 => (x"ff",x"c7",x"49",x"66"),
   753 => (x"87",x"cb",x"02",x"99"),
   754 => (x"1e",x"fa",x"f9",x"c3"),
   755 => (x"d9",x"fc",x"49",x"73"),
   756 => (x"26",x"86",x"c4",x"87"),
   757 => (x"0e",x"87",x"dc",x"f5"),
   758 => (x"5d",x"5c",x"5b",x"5e"),
   759 => (x"d0",x"86",x"f0",x"0e"),
   760 => (x"e4",x"c0",x"59",x"a6"),
   761 => (x"66",x"cc",x"4b",x"66"),
   762 => (x"48",x"87",x"ca",x"02"),
   763 => (x"7e",x"70",x"80",x"c8"),
   764 => (x"c5",x"05",x"bf",x"6e"),
   765 => (x"c3",x"48",x"c0",x"87"),
   766 => (x"66",x"cc",x"87",x"ec"),
   767 => (x"73",x"84",x"d0",x"4c"),
   768 => (x"48",x"a6",x"c4",x"49"),
   769 => (x"66",x"c4",x"78",x"6c"),
   770 => (x"6e",x"80",x"c4",x"81"),
   771 => (x"66",x"c8",x"78",x"bf"),
   772 => (x"87",x"c6",x"06",x"a9"),
   773 => (x"89",x"66",x"c4",x"49"),
   774 => (x"b7",x"c0",x"4b",x"71"),
   775 => (x"87",x"c4",x"01",x"ab"),
   776 => (x"87",x"c2",x"c3",x"48"),
   777 => (x"c7",x"48",x"66",x"c4"),
   778 => (x"7e",x"70",x"98",x"ff"),
   779 => (x"c9",x"c1",x"02",x"6e"),
   780 => (x"49",x"c0",x"c8",x"87"),
   781 => (x"4a",x"71",x"89",x"6e"),
   782 => (x"4d",x"fa",x"f9",x"c3"),
   783 => (x"b7",x"73",x"85",x"6e"),
   784 => (x"87",x"c1",x"06",x"aa"),
   785 => (x"48",x"49",x"72",x"4a"),
   786 => (x"70",x"80",x"66",x"c4"),
   787 => (x"49",x"8b",x"72",x"7c"),
   788 => (x"99",x"71",x"8a",x"c1"),
   789 => (x"c0",x"87",x"d9",x"02"),
   790 => (x"15",x"48",x"66",x"e0"),
   791 => (x"66",x"e0",x"c0",x"50"),
   792 => (x"c0",x"80",x"c1",x"48"),
   793 => (x"72",x"58",x"a6",x"e4"),
   794 => (x"71",x"8a",x"c1",x"49"),
   795 => (x"87",x"e7",x"05",x"99"),
   796 => (x"66",x"d0",x"1e",x"c1"),
   797 => (x"87",x"d1",x"f8",x"49"),
   798 => (x"b7",x"c0",x"86",x"c4"),
   799 => (x"e3",x"c1",x"06",x"ab"),
   800 => (x"66",x"e0",x"c0",x"87"),
   801 => (x"b7",x"ff",x"c7",x"4d"),
   802 => (x"e2",x"c0",x"06",x"ab"),
   803 => (x"d0",x"1e",x"75",x"87"),
   804 => (x"d5",x"f9",x"49",x"66"),
   805 => (x"85",x"c0",x"c8",x"87"),
   806 => (x"c0",x"c8",x"48",x"6c"),
   807 => (x"c8",x"7c",x"70",x"80"),
   808 => (x"1e",x"c1",x"8b",x"c0"),
   809 => (x"f7",x"49",x"66",x"d4"),
   810 => (x"86",x"c8",x"87",x"df"),
   811 => (x"c3",x"87",x"ee",x"c0"),
   812 => (x"d0",x"1e",x"fa",x"f9"),
   813 => (x"f1",x"f8",x"49",x"66"),
   814 => (x"c3",x"86",x"c4",x"87"),
   815 => (x"73",x"4a",x"fa",x"f9"),
   816 => (x"80",x"6c",x"48",x"49"),
   817 => (x"49",x"73",x"7c",x"70"),
   818 => (x"99",x"71",x"8b",x"c1"),
   819 => (x"12",x"87",x"ce",x"02"),
   820 => (x"85",x"c1",x"7d",x"97"),
   821 => (x"8b",x"c1",x"49",x"73"),
   822 => (x"f2",x"05",x"99",x"71"),
   823 => (x"ab",x"b7",x"c0",x"87"),
   824 => (x"87",x"e1",x"fe",x"01"),
   825 => (x"8e",x"f0",x"48",x"c1"),
   826 => (x"0e",x"87",x"c8",x"f1"),
   827 => (x"5d",x"5c",x"5b",x"5e"),
   828 => (x"9b",x"4b",x"71",x"0e"),
   829 => (x"c8",x"87",x"c7",x"02"),
   830 => (x"05",x"6d",x"4d",x"a3"),
   831 => (x"48",x"ff",x"87",x"c5"),
   832 => (x"d0",x"87",x"fd",x"c0"),
   833 => (x"49",x"6c",x"4c",x"a3"),
   834 => (x"05",x"99",x"ff",x"c7"),
   835 => (x"02",x"6c",x"87",x"d8"),
   836 => (x"1e",x"c1",x"87",x"c9"),
   837 => (x"f0",x"f5",x"49",x"73"),
   838 => (x"c3",x"86",x"c4",x"87"),
   839 => (x"73",x"1e",x"fa",x"f9"),
   840 => (x"87",x"c6",x"f7",x"49"),
   841 => (x"4a",x"6c",x"86",x"c4"),
   842 => (x"c4",x"04",x"aa",x"6d"),
   843 => (x"cf",x"48",x"ff",x"87"),
   844 => (x"7c",x"a2",x"c1",x"87"),
   845 => (x"ff",x"c7",x"49",x"72"),
   846 => (x"fa",x"f9",x"c3",x"99"),
   847 => (x"48",x"69",x"97",x"81"),
   848 => (x"1e",x"87",x"f0",x"ef"),
   849 => (x"4b",x"71",x"1e",x"73"),
   850 => (x"e4",x"c0",x"02",x"9b"),
   851 => (x"e7",x"c6",x"c4",x"87"),
   852 => (x"c2",x"4a",x"73",x"5b"),
   853 => (x"fa",x"c1",x"c4",x"8a"),
   854 => (x"c4",x"92",x"49",x"bf"),
   855 => (x"48",x"bf",x"d3",x"c6"),
   856 => (x"c6",x"c4",x"80",x"72"),
   857 => (x"48",x"71",x"58",x"eb"),
   858 => (x"c2",x"c4",x"30",x"c4"),
   859 => (x"ed",x"c0",x"58",x"ca"),
   860 => (x"e3",x"c6",x"c4",x"87"),
   861 => (x"d7",x"c6",x"c4",x"48"),
   862 => (x"c6",x"c4",x"78",x"bf"),
   863 => (x"c6",x"c4",x"48",x"e7"),
   864 => (x"c4",x"78",x"bf",x"db"),
   865 => (x"02",x"bf",x"c2",x"c2"),
   866 => (x"c1",x"c4",x"87",x"c9"),
   867 => (x"c4",x"49",x"bf",x"fa"),
   868 => (x"c4",x"87",x"c7",x"31"),
   869 => (x"49",x"bf",x"df",x"c6"),
   870 => (x"c2",x"c4",x"31",x"c4"),
   871 => (x"d6",x"ee",x"59",x"ca"),
   872 => (x"5b",x"5e",x"0e",x"87"),
   873 => (x"4a",x"71",x"0e",x"5c"),
   874 => (x"9a",x"72",x"4b",x"c0"),
   875 => (x"87",x"e1",x"c0",x"02"),
   876 => (x"9f",x"49",x"a2",x"da"),
   877 => (x"c2",x"c4",x"4b",x"69"),
   878 => (x"cf",x"02",x"bf",x"c2"),
   879 => (x"49",x"a2",x"d4",x"87"),
   880 => (x"4c",x"49",x"69",x"9f"),
   881 => (x"9c",x"ff",x"ff",x"c0"),
   882 => (x"87",x"c2",x"34",x"d0"),
   883 => (x"49",x"74",x"4c",x"c0"),
   884 => (x"fd",x"49",x"73",x"b3"),
   885 => (x"dc",x"ed",x"87",x"ed"),
   886 => (x"5b",x"5e",x"0e",x"87"),
   887 => (x"f4",x"0e",x"5d",x"5c"),
   888 => (x"c0",x"4a",x"71",x"86"),
   889 => (x"02",x"9a",x"72",x"7e"),
   890 => (x"f9",x"c3",x"87",x"d8"),
   891 => (x"78",x"c0",x"48",x"f6"),
   892 => (x"48",x"ee",x"f9",x"c3"),
   893 => (x"bf",x"e7",x"c6",x"c4"),
   894 => (x"f2",x"f9",x"c3",x"78"),
   895 => (x"e3",x"c6",x"c4",x"48"),
   896 => (x"c2",x"c4",x"78",x"bf"),
   897 => (x"50",x"c0",x"48",x"d7"),
   898 => (x"bf",x"c6",x"c2",x"c4"),
   899 => (x"f6",x"f9",x"c3",x"49"),
   900 => (x"aa",x"71",x"4a",x"bf"),
   901 => (x"87",x"c0",x"c4",x"03"),
   902 => (x"99",x"cf",x"49",x"72"),
   903 => (x"87",x"e1",x"c0",x"05"),
   904 => (x"1e",x"fa",x"f9",x"c3"),
   905 => (x"bf",x"ee",x"f9",x"c3"),
   906 => (x"ee",x"f9",x"c3",x"49"),
   907 => (x"78",x"a1",x"c1",x"48"),
   908 => (x"c0",x"de",x"ff",x"71"),
   909 => (x"c0",x"86",x"c4",x"87"),
   910 => (x"c3",x"48",x"ed",x"fe"),
   911 => (x"cc",x"78",x"fa",x"f9"),
   912 => (x"ed",x"fe",x"c0",x"87"),
   913 => (x"e0",x"c0",x"48",x"bf"),
   914 => (x"f1",x"fe",x"c0",x"80"),
   915 => (x"f6",x"f9",x"c3",x"58"),
   916 => (x"80",x"c1",x"48",x"bf"),
   917 => (x"58",x"fa",x"f9",x"c3"),
   918 => (x"00",x"0f",x"ad",x"27"),
   919 => (x"bf",x"97",x"bf",x"00"),
   920 => (x"c2",x"02",x"9d",x"4d"),
   921 => (x"e5",x"c3",x"87",x"e2"),
   922 => (x"db",x"c2",x"02",x"ad"),
   923 => (x"ed",x"fe",x"c0",x"87"),
   924 => (x"a3",x"cb",x"4b",x"bf"),
   925 => (x"cf",x"4c",x"11",x"49"),
   926 => (x"d2",x"c1",x"05",x"ac"),
   927 => (x"df",x"49",x"75",x"87"),
   928 => (x"cd",x"89",x"c1",x"99"),
   929 => (x"ca",x"c2",x"c4",x"91"),
   930 => (x"4a",x"a3",x"c1",x"81"),
   931 => (x"a3",x"c3",x"51",x"12"),
   932 => (x"c5",x"51",x"12",x"4a"),
   933 => (x"51",x"12",x"4a",x"a3"),
   934 => (x"12",x"4a",x"a3",x"c7"),
   935 => (x"4a",x"a3",x"c9",x"51"),
   936 => (x"a3",x"ce",x"51",x"12"),
   937 => (x"d0",x"51",x"12",x"4a"),
   938 => (x"51",x"12",x"4a",x"a3"),
   939 => (x"12",x"4a",x"a3",x"d2"),
   940 => (x"4a",x"a3",x"d4",x"51"),
   941 => (x"a3",x"d6",x"51",x"12"),
   942 => (x"d8",x"51",x"12",x"4a"),
   943 => (x"51",x"12",x"4a",x"a3"),
   944 => (x"12",x"4a",x"a3",x"dc"),
   945 => (x"4a",x"a3",x"de",x"51"),
   946 => (x"7e",x"c1",x"51",x"12"),
   947 => (x"74",x"87",x"f9",x"c0"),
   948 => (x"05",x"99",x"c8",x"49"),
   949 => (x"74",x"87",x"ea",x"c0"),
   950 => (x"05",x"99",x"d0",x"49"),
   951 => (x"66",x"dc",x"87",x"d0"),
   952 => (x"87",x"ca",x"c0",x"02"),
   953 => (x"66",x"dc",x"49",x"73"),
   954 => (x"02",x"98",x"70",x"0f"),
   955 => (x"05",x"6e",x"87",x"d3"),
   956 => (x"c4",x"87",x"c6",x"c0"),
   957 => (x"c0",x"48",x"ca",x"c2"),
   958 => (x"ed",x"fe",x"c0",x"50"),
   959 => (x"e7",x"c2",x"48",x"bf"),
   960 => (x"d7",x"c2",x"c4",x"87"),
   961 => (x"7e",x"50",x"c0",x"48"),
   962 => (x"bf",x"c6",x"c2",x"c4"),
   963 => (x"f6",x"f9",x"c3",x"49"),
   964 => (x"aa",x"71",x"4a",x"bf"),
   965 => (x"87",x"c0",x"fc",x"04"),
   966 => (x"bf",x"e7",x"c6",x"c4"),
   967 => (x"87",x"c8",x"c0",x"05"),
   968 => (x"bf",x"c2",x"c2",x"c4"),
   969 => (x"87",x"fe",x"c1",x"02"),
   970 => (x"48",x"f1",x"fe",x"c0"),
   971 => (x"f9",x"c3",x"78",x"ff"),
   972 => (x"e8",x"49",x"bf",x"f2"),
   973 => (x"49",x"70",x"87",x"c5"),
   974 => (x"59",x"f6",x"f9",x"c3"),
   975 => (x"c3",x"48",x"a6",x"c4"),
   976 => (x"78",x"bf",x"f2",x"f9"),
   977 => (x"bf",x"c2",x"c2",x"c4"),
   978 => (x"87",x"d8",x"c0",x"02"),
   979 => (x"cf",x"49",x"66",x"c4"),
   980 => (x"f8",x"ff",x"ff",x"ff"),
   981 => (x"c0",x"02",x"a9",x"99"),
   982 => (x"4d",x"c0",x"87",x"c5"),
   983 => (x"c1",x"87",x"e1",x"c0"),
   984 => (x"87",x"dc",x"c0",x"4d"),
   985 => (x"cf",x"49",x"66",x"c4"),
   986 => (x"a9",x"99",x"f8",x"ff"),
   987 => (x"87",x"c8",x"c0",x"02"),
   988 => (x"c0",x"48",x"a6",x"c8"),
   989 => (x"87",x"c5",x"c0",x"78"),
   990 => (x"c1",x"48",x"a6",x"c8"),
   991 => (x"4d",x"66",x"c8",x"78"),
   992 => (x"c0",x"05",x"9d",x"75"),
   993 => (x"66",x"c4",x"87",x"e0"),
   994 => (x"c4",x"89",x"c2",x"49"),
   995 => (x"4a",x"bf",x"fa",x"c1"),
   996 => (x"d3",x"c6",x"c4",x"91"),
   997 => (x"f9",x"c3",x"4a",x"bf"),
   998 => (x"a1",x"72",x"48",x"ee"),
   999 => (x"f6",x"f9",x"c3",x"78"),
  1000 => (x"f9",x"78",x"c0",x"48"),
  1001 => (x"48",x"c0",x"87",x"e2"),
  1002 => (x"c6",x"e6",x"8e",x"f4"),
  1003 => (x"00",x"00",x"00",x"87"),
  1004 => (x"ff",x"ff",x"ff",x"00"),
  1005 => (x"00",x"0f",x"bd",x"ff"),
  1006 => (x"00",x"0f",x"c6",x"00"),
  1007 => (x"54",x"41",x"46",x"00"),
  1008 => (x"20",x"20",x"32",x"33"),
  1009 => (x"41",x"46",x"00",x"20"),
  1010 => (x"20",x"36",x"31",x"54"),
  1011 => (x"1e",x"00",x"20",x"20"),
  1012 => (x"c3",x"48",x"d4",x"ff"),
  1013 => (x"48",x"68",x"78",x"ff"),
  1014 => (x"ff",x"1e",x"4f",x"26"),
  1015 => (x"ff",x"c3",x"48",x"d4"),
  1016 => (x"48",x"d0",x"ff",x"78"),
  1017 => (x"ff",x"78",x"e1",x"c8"),
  1018 => (x"78",x"d4",x"48",x"d4"),
  1019 => (x"48",x"eb",x"c6",x"c4"),
  1020 => (x"50",x"bf",x"d4",x"ff"),
  1021 => (x"ff",x"1e",x"4f",x"26"),
  1022 => (x"e0",x"c0",x"48",x"d0"),
  1023 => (x"1e",x"4f",x"26",x"78"),
  1024 => (x"70",x"87",x"cc",x"ff"),
  1025 => (x"c6",x"02",x"99",x"49"),
  1026 => (x"a9",x"fb",x"c0",x"87"),
  1027 => (x"71",x"87",x"f1",x"05"),
  1028 => (x"0e",x"4f",x"26",x"48"),
  1029 => (x"0e",x"5c",x"5b",x"5e"),
  1030 => (x"4c",x"c0",x"4b",x"71"),
  1031 => (x"70",x"87",x"f0",x"fe"),
  1032 => (x"c0",x"02",x"99",x"49"),
  1033 => (x"ec",x"c0",x"87",x"f9"),
  1034 => (x"f2",x"c0",x"02",x"a9"),
  1035 => (x"a9",x"fb",x"c0",x"87"),
  1036 => (x"87",x"eb",x"c0",x"02"),
  1037 => (x"ac",x"b7",x"66",x"cc"),
  1038 => (x"d0",x"87",x"c7",x"03"),
  1039 => (x"87",x"c2",x"02",x"66"),
  1040 => (x"99",x"71",x"53",x"71"),
  1041 => (x"c1",x"87",x"c2",x"02"),
  1042 => (x"87",x"c3",x"fe",x"84"),
  1043 => (x"02",x"99",x"49",x"70"),
  1044 => (x"ec",x"c0",x"87",x"cd"),
  1045 => (x"87",x"c7",x"02",x"a9"),
  1046 => (x"05",x"a9",x"fb",x"c0"),
  1047 => (x"d0",x"87",x"d5",x"ff"),
  1048 => (x"87",x"c3",x"02",x"66"),
  1049 => (x"c0",x"7b",x"97",x"c0"),
  1050 => (x"c4",x"05",x"a9",x"ec"),
  1051 => (x"c5",x"4a",x"74",x"87"),
  1052 => (x"c0",x"4a",x"74",x"87"),
  1053 => (x"48",x"72",x"8a",x"0a"),
  1054 => (x"4d",x"26",x"87",x"c2"),
  1055 => (x"4b",x"26",x"4c",x"26"),
  1056 => (x"fd",x"1e",x"4f",x"26"),
  1057 => (x"49",x"70",x"87",x"c9"),
  1058 => (x"a9",x"b7",x"f0",x"c0"),
  1059 => (x"c0",x"87",x"ca",x"04"),
  1060 => (x"01",x"a9",x"b7",x"f9"),
  1061 => (x"f0",x"c0",x"87",x"c3"),
  1062 => (x"b7",x"c1",x"c1",x"89"),
  1063 => (x"87",x"ca",x"04",x"a9"),
  1064 => (x"a9",x"b7",x"da",x"c1"),
  1065 => (x"c0",x"87",x"c3",x"01"),
  1066 => (x"48",x"71",x"89",x"f7"),
  1067 => (x"5e",x"0e",x"4f",x"26"),
  1068 => (x"71",x"0e",x"5c",x"5b"),
  1069 => (x"4c",x"d4",x"ff",x"4a"),
  1070 => (x"ea",x"c0",x"49",x"72"),
  1071 => (x"9b",x"4b",x"70",x"87"),
  1072 => (x"c1",x"87",x"c2",x"02"),
  1073 => (x"48",x"d0",x"ff",x"8b"),
  1074 => (x"c1",x"78",x"c5",x"c8"),
  1075 => (x"49",x"73",x"7c",x"d5"),
  1076 => (x"f7",x"c3",x"31",x"c6"),
  1077 => (x"4a",x"bf",x"97",x"eb"),
  1078 => (x"70",x"b0",x"71",x"48"),
  1079 => (x"48",x"d0",x"ff",x"7c"),
  1080 => (x"48",x"73",x"78",x"c4"),
  1081 => (x"0e",x"87",x"d5",x"fe"),
  1082 => (x"5d",x"5c",x"5b",x"5e"),
  1083 => (x"71",x"86",x"f8",x"0e"),
  1084 => (x"fb",x"7e",x"c0",x"4c"),
  1085 => (x"4b",x"c0",x"87",x"e4"),
  1086 => (x"97",x"d4",x"c6",x"c1"),
  1087 => (x"a9",x"c0",x"49",x"bf"),
  1088 => (x"fb",x"87",x"cf",x"04"),
  1089 => (x"83",x"c1",x"87",x"f9"),
  1090 => (x"97",x"d4",x"c6",x"c1"),
  1091 => (x"06",x"ab",x"49",x"bf"),
  1092 => (x"c6",x"c1",x"87",x"f1"),
  1093 => (x"02",x"bf",x"97",x"d4"),
  1094 => (x"f2",x"fa",x"87",x"cf"),
  1095 => (x"99",x"49",x"70",x"87"),
  1096 => (x"c0",x"87",x"c6",x"02"),
  1097 => (x"f1",x"05",x"a9",x"ec"),
  1098 => (x"fa",x"4b",x"c0",x"87"),
  1099 => (x"4d",x"70",x"87",x"e1"),
  1100 => (x"c8",x"87",x"dc",x"fa"),
  1101 => (x"d6",x"fa",x"58",x"a6"),
  1102 => (x"c1",x"4a",x"70",x"87"),
  1103 => (x"49",x"a4",x"c8",x"83"),
  1104 => (x"ad",x"49",x"69",x"97"),
  1105 => (x"c0",x"87",x"c7",x"02"),
  1106 => (x"c0",x"05",x"ad",x"ff"),
  1107 => (x"a4",x"c9",x"87",x"e7"),
  1108 => (x"49",x"69",x"97",x"49"),
  1109 => (x"02",x"a9",x"66",x"c4"),
  1110 => (x"c0",x"48",x"87",x"c7"),
  1111 => (x"d4",x"05",x"a8",x"ff"),
  1112 => (x"49",x"a4",x"ca",x"87"),
  1113 => (x"aa",x"49",x"69",x"97"),
  1114 => (x"c0",x"87",x"c6",x"02"),
  1115 => (x"c4",x"05",x"aa",x"ff"),
  1116 => (x"d0",x"7e",x"c1",x"87"),
  1117 => (x"ad",x"ec",x"c0",x"87"),
  1118 => (x"c0",x"87",x"c6",x"02"),
  1119 => (x"c4",x"05",x"ad",x"fb"),
  1120 => (x"c1",x"4b",x"c0",x"87"),
  1121 => (x"fe",x"02",x"6e",x"7e"),
  1122 => (x"e9",x"f9",x"87",x"e1"),
  1123 => (x"f8",x"48",x"73",x"87"),
  1124 => (x"87",x"e6",x"fb",x"8e"),
  1125 => (x"5b",x"5e",x"0e",x"00"),
  1126 => (x"1e",x"0e",x"5d",x"5c"),
  1127 => (x"4c",x"c0",x"4b",x"71"),
  1128 => (x"c0",x"04",x"ab",x"4d"),
  1129 => (x"c3",x"c1",x"87",x"e8"),
  1130 => (x"9d",x"75",x"1e",x"e7"),
  1131 => (x"c0",x"87",x"c4",x"02"),
  1132 => (x"c1",x"87",x"c2",x"4a"),
  1133 => (x"f0",x"49",x"72",x"4a"),
  1134 => (x"86",x"c4",x"87",x"df"),
  1135 => (x"84",x"c1",x"7e",x"70"),
  1136 => (x"87",x"c2",x"05",x"6e"),
  1137 => (x"85",x"c1",x"4c",x"73"),
  1138 => (x"ff",x"06",x"ac",x"73"),
  1139 => (x"48",x"6e",x"87",x"d8"),
  1140 => (x"26",x"4d",x"26",x"26"),
  1141 => (x"26",x"4b",x"26",x"4c"),
  1142 => (x"4a",x"71",x"1e",x"4f"),
  1143 => (x"99",x"ff",x"c3",x"49"),
  1144 => (x"71",x"48",x"d4",x"ff"),
  1145 => (x"c8",x"49",x"72",x"78"),
  1146 => (x"ff",x"c3",x"29",x"b7"),
  1147 => (x"72",x"78",x"71",x"99"),
  1148 => (x"29",x"b7",x"d0",x"49"),
  1149 => (x"71",x"99",x"ff",x"c3"),
  1150 => (x"d8",x"49",x"72",x"78"),
  1151 => (x"ff",x"c3",x"29",x"b7"),
  1152 => (x"26",x"78",x"71",x"99"),
  1153 => (x"5b",x"5e",x"0e",x"4f"),
  1154 => (x"1e",x"0e",x"5d",x"5c"),
  1155 => (x"4b",x"c0",x"4a",x"71"),
  1156 => (x"e3",x"c1",x"49",x"72"),
  1157 => (x"98",x"70",x"87",x"c5"),
  1158 => (x"c1",x"87",x"da",x"05"),
  1159 => (x"c1",x"49",x"74",x"4c"),
  1160 => (x"70",x"87",x"d2",x"e4"),
  1161 => (x"87",x"c2",x"05",x"98"),
  1162 => (x"84",x"c1",x"4b",x"c1"),
  1163 => (x"bf",x"ce",x"cb",x"c4"),
  1164 => (x"e8",x"06",x"ac",x"b7"),
  1165 => (x"48",x"d0",x"ff",x"87"),
  1166 => (x"ff",x"78",x"e1",x"c8"),
  1167 => (x"78",x"dd",x"48",x"d4"),
  1168 => (x"c7",x"02",x"9b",x"73"),
  1169 => (x"f6",x"cb",x"c4",x"87"),
  1170 => (x"87",x"c2",x"4d",x"bf"),
  1171 => (x"49",x"75",x"4d",x"c0"),
  1172 => (x"73",x"87",x"c6",x"fe"),
  1173 => (x"87",x"c7",x"02",x"9b"),
  1174 => (x"bf",x"f6",x"cb",x"c4"),
  1175 => (x"c0",x"87",x"c2",x"7e"),
  1176 => (x"fd",x"49",x"6e",x"7e"),
  1177 => (x"49",x"c0",x"87",x"f3"),
  1178 => (x"c0",x"87",x"ee",x"fd"),
  1179 => (x"87",x"e9",x"fd",x"49"),
  1180 => (x"c0",x"48",x"d0",x"ff"),
  1181 => (x"1e",x"c1",x"78",x"e0"),
  1182 => (x"f2",x"c0",x"49",x"dc"),
  1183 => (x"48",x"73",x"87",x"ca"),
  1184 => (x"cc",x"fd",x"8e",x"f8"),
  1185 => (x"5b",x"5e",x"0e",x"87"),
  1186 => (x"1e",x"0e",x"5d",x"5c"),
  1187 => (x"de",x"49",x"4c",x"71"),
  1188 => (x"c5",x"c7",x"c4",x"91"),
  1189 => (x"97",x"85",x"71",x"4d"),
  1190 => (x"dd",x"c1",x"02",x"6d"),
  1191 => (x"f0",x"c6",x"c4",x"87"),
  1192 => (x"82",x"74",x"4a",x"bf"),
  1193 => (x"ec",x"fb",x"49",x"72"),
  1194 => (x"6e",x"7e",x"70",x"87"),
  1195 => (x"87",x"f3",x"c0",x"02"),
  1196 => (x"4b",x"f8",x"c6",x"c4"),
  1197 => (x"49",x"cb",x"4a",x"6e"),
  1198 => (x"87",x"fd",x"f7",x"fe"),
  1199 => (x"93",x"cb",x"4b",x"74"),
  1200 => (x"83",x"d3",x"ed",x"c1"),
  1201 => (x"cb",x"c1",x"83",x"c4"),
  1202 => (x"49",x"74",x"7b",x"fe"),
  1203 => (x"87",x"ee",x"c4",x"c1"),
  1204 => (x"c7",x"c4",x"7b",x"75"),
  1205 => (x"49",x"bf",x"97",x"c4"),
  1206 => (x"f8",x"c6",x"c4",x"1e"),
  1207 => (x"ff",x"ea",x"c2",x"49"),
  1208 => (x"74",x"86",x"c4",x"87"),
  1209 => (x"d5",x"c4",x"c1",x"49"),
  1210 => (x"c1",x"49",x"c0",x"87"),
  1211 => (x"c4",x"87",x"f4",x"c5"),
  1212 => (x"c0",x"48",x"ec",x"c6"),
  1213 => (x"dd",x"49",x"c1",x"78"),
  1214 => (x"fb",x"26",x"87",x"c1"),
  1215 => (x"6f",x"4c",x"87",x"d3"),
  1216 => (x"6e",x"69",x"64",x"61"),
  1217 => (x"2e",x"2e",x"2e",x"67"),
  1218 => (x"5b",x"5e",x"0e",x"00"),
  1219 => (x"4b",x"71",x"0e",x"5c"),
  1220 => (x"f0",x"c6",x"c4",x"4a"),
  1221 => (x"49",x"72",x"82",x"bf"),
  1222 => (x"70",x"87",x"fa",x"f9"),
  1223 => (x"c4",x"02",x"9c",x"4c"),
  1224 => (x"fc",x"e9",x"49",x"87"),
  1225 => (x"f0",x"c6",x"c4",x"87"),
  1226 => (x"c1",x"78",x"c0",x"48"),
  1227 => (x"87",x"cb",x"dc",x"49"),
  1228 => (x"0e",x"87",x"e0",x"fa"),
  1229 => (x"5d",x"5c",x"5b",x"5e"),
  1230 => (x"c3",x"86",x"f4",x"0e"),
  1231 => (x"c0",x"4d",x"fa",x"f9"),
  1232 => (x"48",x"a6",x"c4",x"4c"),
  1233 => (x"c6",x"c4",x"78",x"c0"),
  1234 => (x"c0",x"49",x"bf",x"f0"),
  1235 => (x"c1",x"c1",x"06",x"a9"),
  1236 => (x"fa",x"f9",x"c3",x"87"),
  1237 => (x"c0",x"02",x"98",x"48"),
  1238 => (x"c3",x"c1",x"87",x"f8"),
  1239 => (x"66",x"c8",x"1e",x"e7"),
  1240 => (x"c4",x"87",x"c7",x"02"),
  1241 => (x"78",x"c0",x"48",x"a6"),
  1242 => (x"a6",x"c4",x"87",x"c5"),
  1243 => (x"c4",x"78",x"c1",x"48"),
  1244 => (x"e4",x"e9",x"49",x"66"),
  1245 => (x"70",x"86",x"c4",x"87"),
  1246 => (x"c4",x"84",x"c1",x"4d"),
  1247 => (x"80",x"c1",x"48",x"66"),
  1248 => (x"c4",x"58",x"a6",x"c8"),
  1249 => (x"49",x"bf",x"f0",x"c6"),
  1250 => (x"87",x"c6",x"03",x"ac"),
  1251 => (x"ff",x"05",x"9d",x"75"),
  1252 => (x"4c",x"c0",x"87",x"c8"),
  1253 => (x"c3",x"02",x"9d",x"75"),
  1254 => (x"c3",x"c1",x"87",x"e0"),
  1255 => (x"66",x"c8",x"1e",x"e7"),
  1256 => (x"cc",x"87",x"c7",x"02"),
  1257 => (x"78",x"c0",x"48",x"a6"),
  1258 => (x"a6",x"cc",x"87",x"c5"),
  1259 => (x"cc",x"78",x"c1",x"48"),
  1260 => (x"e4",x"e8",x"49",x"66"),
  1261 => (x"70",x"86",x"c4",x"87"),
  1262 => (x"c2",x"02",x"6e",x"7e"),
  1263 => (x"49",x"6e",x"87",x"e9"),
  1264 => (x"69",x"97",x"81",x"cb"),
  1265 => (x"02",x"99",x"d0",x"49"),
  1266 => (x"c1",x"87",x"d6",x"c1"),
  1267 => (x"74",x"4a",x"c9",x"cc"),
  1268 => (x"c1",x"91",x"cb",x"49"),
  1269 => (x"72",x"81",x"d3",x"ed"),
  1270 => (x"c3",x"81",x"c8",x"79"),
  1271 => (x"49",x"74",x"51",x"ff"),
  1272 => (x"c7",x"c4",x"91",x"de"),
  1273 => (x"85",x"71",x"4d",x"c5"),
  1274 => (x"7d",x"97",x"c1",x"c2"),
  1275 => (x"c0",x"49",x"a5",x"c1"),
  1276 => (x"c2",x"c4",x"51",x"e0"),
  1277 => (x"02",x"bf",x"97",x"ca"),
  1278 => (x"84",x"c1",x"87",x"d2"),
  1279 => (x"c4",x"4b",x"a5",x"c2"),
  1280 => (x"db",x"4a",x"ca",x"c2"),
  1281 => (x"f0",x"f2",x"fe",x"49"),
  1282 => (x"87",x"db",x"c1",x"87"),
  1283 => (x"c0",x"49",x"a5",x"cd"),
  1284 => (x"c2",x"84",x"c1",x"51"),
  1285 => (x"4a",x"6e",x"4b",x"a5"),
  1286 => (x"f2",x"fe",x"49",x"cb"),
  1287 => (x"c6",x"c1",x"87",x"db"),
  1288 => (x"c5",x"ca",x"c1",x"87"),
  1289 => (x"cb",x"49",x"74",x"4a"),
  1290 => (x"d3",x"ed",x"c1",x"91"),
  1291 => (x"c4",x"79",x"72",x"81"),
  1292 => (x"bf",x"97",x"ca",x"c2"),
  1293 => (x"74",x"87",x"d8",x"02"),
  1294 => (x"c1",x"91",x"de",x"49"),
  1295 => (x"c5",x"c7",x"c4",x"84"),
  1296 => (x"c4",x"83",x"71",x"4b"),
  1297 => (x"dd",x"4a",x"ca",x"c2"),
  1298 => (x"ec",x"f1",x"fe",x"49"),
  1299 => (x"74",x"87",x"d8",x"87"),
  1300 => (x"c4",x"93",x"de",x"4b"),
  1301 => (x"cb",x"83",x"c5",x"c7"),
  1302 => (x"51",x"c0",x"49",x"a3"),
  1303 => (x"6e",x"73",x"84",x"c1"),
  1304 => (x"fe",x"49",x"cb",x"4a"),
  1305 => (x"c4",x"87",x"d2",x"f1"),
  1306 => (x"80",x"c1",x"48",x"66"),
  1307 => (x"c7",x"58",x"a6",x"c8"),
  1308 => (x"c5",x"c0",x"03",x"ac"),
  1309 => (x"fc",x"05",x"6e",x"87"),
  1310 => (x"48",x"74",x"87",x"e0"),
  1311 => (x"d0",x"f5",x"8e",x"f4"),
  1312 => (x"1e",x"73",x"1e",x"87"),
  1313 => (x"cb",x"49",x"4b",x"71"),
  1314 => (x"d3",x"ed",x"c1",x"91"),
  1315 => (x"4a",x"a1",x"c8",x"81"),
  1316 => (x"48",x"eb",x"f7",x"c3"),
  1317 => (x"a1",x"c9",x"50",x"12"),
  1318 => (x"d4",x"c6",x"c1",x"4a"),
  1319 => (x"ca",x"50",x"12",x"48"),
  1320 => (x"c4",x"c7",x"c4",x"81"),
  1321 => (x"c4",x"50",x"11",x"48"),
  1322 => (x"bf",x"97",x"c4",x"c7"),
  1323 => (x"49",x"c0",x"1e",x"49"),
  1324 => (x"87",x"ec",x"e3",x"c2"),
  1325 => (x"48",x"ec",x"c6",x"c4"),
  1326 => (x"49",x"c1",x"78",x"de"),
  1327 => (x"26",x"87",x"fc",x"d5"),
  1328 => (x"1e",x"87",x"d2",x"f4"),
  1329 => (x"cb",x"49",x"4a",x"71"),
  1330 => (x"d3",x"ed",x"c1",x"91"),
  1331 => (x"11",x"81",x"c8",x"81"),
  1332 => (x"f0",x"c6",x"c4",x"48"),
  1333 => (x"f0",x"c6",x"c4",x"58"),
  1334 => (x"c1",x"78",x"c0",x"48"),
  1335 => (x"87",x"db",x"d5",x"49"),
  1336 => (x"c0",x"1e",x"4f",x"26"),
  1337 => (x"fa",x"fd",x"c0",x"49"),
  1338 => (x"1e",x"4f",x"26",x"87"),
  1339 => (x"d2",x"02",x"99",x"71"),
  1340 => (x"e8",x"ee",x"c1",x"87"),
  1341 => (x"f7",x"50",x"c0",x"48"),
  1342 => (x"c3",x"d3",x"c1",x"80"),
  1343 => (x"cc",x"ed",x"c1",x"40"),
  1344 => (x"c1",x"87",x"ce",x"78"),
  1345 => (x"c1",x"48",x"e4",x"ee"),
  1346 => (x"fc",x"78",x"c5",x"ed"),
  1347 => (x"e2",x"d3",x"c1",x"80"),
  1348 => (x"0e",x"4f",x"26",x"78"),
  1349 => (x"0e",x"5c",x"5b",x"5e"),
  1350 => (x"cb",x"4a",x"4c",x"71"),
  1351 => (x"d3",x"ed",x"c1",x"92"),
  1352 => (x"49",x"a2",x"c8",x"82"),
  1353 => (x"97",x"4b",x"a2",x"c9"),
  1354 => (x"97",x"1e",x"4b",x"6b"),
  1355 => (x"ca",x"1e",x"49",x"69"),
  1356 => (x"c0",x"49",x"12",x"82"),
  1357 => (x"c0",x"87",x"f5",x"e8"),
  1358 => (x"87",x"ff",x"d3",x"49"),
  1359 => (x"fa",x"c0",x"49",x"74"),
  1360 => (x"8e",x"f8",x"87",x"fc"),
  1361 => (x"1e",x"87",x"cc",x"f2"),
  1362 => (x"4b",x"71",x"1e",x"73"),
  1363 => (x"87",x"c3",x"ff",x"49"),
  1364 => (x"fe",x"fe",x"49",x"73"),
  1365 => (x"87",x"fd",x"f1",x"87"),
  1366 => (x"71",x"1e",x"73",x"1e"),
  1367 => (x"4a",x"a3",x"c6",x"4b"),
  1368 => (x"c1",x"87",x"db",x"02"),
  1369 => (x"87",x"d6",x"02",x"8a"),
  1370 => (x"da",x"c1",x"02",x"8a"),
  1371 => (x"c0",x"02",x"8a",x"87"),
  1372 => (x"02",x"8a",x"87",x"fc"),
  1373 => (x"8a",x"87",x"e1",x"c0"),
  1374 => (x"c1",x"87",x"cb",x"02"),
  1375 => (x"49",x"c7",x"87",x"db"),
  1376 => (x"c1",x"87",x"c0",x"fd"),
  1377 => (x"c6",x"c4",x"87",x"de"),
  1378 => (x"c1",x"02",x"bf",x"f0"),
  1379 => (x"c1",x"48",x"87",x"cb"),
  1380 => (x"f4",x"c6",x"c4",x"88"),
  1381 => (x"87",x"c1",x"c1",x"58"),
  1382 => (x"bf",x"f4",x"c6",x"c4"),
  1383 => (x"87",x"f9",x"c0",x"02"),
  1384 => (x"bf",x"f0",x"c6",x"c4"),
  1385 => (x"c4",x"80",x"c1",x"48"),
  1386 => (x"c0",x"58",x"f4",x"c6"),
  1387 => (x"c6",x"c4",x"87",x"eb"),
  1388 => (x"c6",x"49",x"bf",x"f0"),
  1389 => (x"f4",x"c6",x"c4",x"89"),
  1390 => (x"a9",x"b7",x"c0",x"59"),
  1391 => (x"c4",x"87",x"da",x"03"),
  1392 => (x"c0",x"48",x"f0",x"c6"),
  1393 => (x"c4",x"87",x"d2",x"78"),
  1394 => (x"02",x"bf",x"f4",x"c6"),
  1395 => (x"c6",x"c4",x"87",x"cb"),
  1396 => (x"c6",x"48",x"bf",x"f0"),
  1397 => (x"f4",x"c6",x"c4",x"80"),
  1398 => (x"d1",x"49",x"c0",x"58"),
  1399 => (x"49",x"73",x"87",x"dd"),
  1400 => (x"87",x"da",x"f8",x"c0"),
  1401 => (x"0e",x"87",x"ee",x"ef"),
  1402 => (x"0e",x"5c",x"5b",x"5e"),
  1403 => (x"66",x"cc",x"4c",x"71"),
  1404 => (x"cb",x"4b",x"74",x"1e"),
  1405 => (x"d3",x"ed",x"c1",x"93"),
  1406 => (x"4a",x"a3",x"c4",x"83"),
  1407 => (x"eb",x"fe",x"49",x"6a"),
  1408 => (x"d2",x"c1",x"87",x"c7"),
  1409 => (x"a3",x"c8",x"7b",x"c1"),
  1410 => (x"51",x"66",x"d4",x"49"),
  1411 => (x"d8",x"49",x"a3",x"c9"),
  1412 => (x"a3",x"ca",x"51",x"66"),
  1413 => (x"51",x"66",x"dc",x"49"),
  1414 => (x"87",x"f7",x"ee",x"26"),
  1415 => (x"5c",x"5b",x"5e",x"0e"),
  1416 => (x"d0",x"ff",x"0e",x"5d"),
  1417 => (x"59",x"a6",x"d8",x"86"),
  1418 => (x"c0",x"48",x"a6",x"c4"),
  1419 => (x"c1",x"80",x"c4",x"78"),
  1420 => (x"c4",x"78",x"66",x"c4"),
  1421 => (x"c4",x"78",x"c1",x"80"),
  1422 => (x"c4",x"78",x"c1",x"80"),
  1423 => (x"c1",x"48",x"f4",x"c6"),
  1424 => (x"ec",x"c6",x"c4",x"78"),
  1425 => (x"a8",x"de",x"48",x"bf"),
  1426 => (x"f3",x"87",x"cb",x"05"),
  1427 => (x"49",x"70",x"87",x"e5"),
  1428 => (x"ce",x"59",x"a6",x"c8"),
  1429 => (x"c1",x"e6",x"87",x"ed"),
  1430 => (x"87",x"e3",x"e6",x"87"),
  1431 => (x"70",x"87",x"f0",x"e5"),
  1432 => (x"ac",x"fb",x"c0",x"4c"),
  1433 => (x"87",x"d0",x"c1",x"02"),
  1434 => (x"c1",x"05",x"66",x"d4"),
  1435 => (x"1e",x"c0",x"87",x"c2"),
  1436 => (x"c1",x"1e",x"c1",x"1e"),
  1437 => (x"c0",x"1e",x"c6",x"ef"),
  1438 => (x"87",x"eb",x"fd",x"49"),
  1439 => (x"4a",x"66",x"d0",x"c1"),
  1440 => (x"49",x"6a",x"82",x"c4"),
  1441 => (x"51",x"74",x"81",x"c7"),
  1442 => (x"1e",x"d8",x"1e",x"c1"),
  1443 => (x"81",x"c8",x"49",x"6a"),
  1444 => (x"d8",x"87",x"c0",x"e6"),
  1445 => (x"66",x"c4",x"c1",x"86"),
  1446 => (x"01",x"a8",x"c0",x"48"),
  1447 => (x"a6",x"c4",x"87",x"c7"),
  1448 => (x"ce",x"78",x"c1",x"48"),
  1449 => (x"66",x"c4",x"c1",x"87"),
  1450 => (x"cc",x"88",x"c1",x"48"),
  1451 => (x"87",x"c3",x"58",x"a6"),
  1452 => (x"cc",x"87",x"cc",x"e5"),
  1453 => (x"78",x"c2",x"48",x"a6"),
  1454 => (x"cd",x"02",x"9c",x"74"),
  1455 => (x"66",x"c4",x"87",x"c1"),
  1456 => (x"66",x"c8",x"c1",x"48"),
  1457 => (x"f6",x"cc",x"03",x"a8"),
  1458 => (x"48",x"a6",x"d8",x"87"),
  1459 => (x"80",x"c4",x"78",x"c0"),
  1460 => (x"fa",x"e3",x"78",x"c0"),
  1461 => (x"c1",x"4c",x"70",x"87"),
  1462 => (x"c2",x"05",x"ac",x"d0"),
  1463 => (x"66",x"dc",x"87",x"d7"),
  1464 => (x"87",x"de",x"e6",x"7e"),
  1465 => (x"e0",x"c0",x"49",x"70"),
  1466 => (x"e2",x"e3",x"59",x"a6"),
  1467 => (x"c0",x"4c",x"70",x"87"),
  1468 => (x"c1",x"05",x"ac",x"ec"),
  1469 => (x"66",x"c4",x"87",x"ea"),
  1470 => (x"c1",x"91",x"cb",x"49"),
  1471 => (x"c4",x"81",x"66",x"c0"),
  1472 => (x"4d",x"6a",x"4a",x"a1"),
  1473 => (x"dc",x"4a",x"a1",x"c8"),
  1474 => (x"d3",x"c1",x"52",x"66"),
  1475 => (x"fe",x"e2",x"79",x"c3"),
  1476 => (x"9c",x"4c",x"70",x"87"),
  1477 => (x"c0",x"87",x"d8",x"02"),
  1478 => (x"d2",x"02",x"ac",x"fb"),
  1479 => (x"e2",x"55",x"74",x"87"),
  1480 => (x"4c",x"70",x"87",x"ed"),
  1481 => (x"87",x"c7",x"02",x"9c"),
  1482 => (x"05",x"ac",x"fb",x"c0"),
  1483 => (x"c0",x"87",x"ee",x"ff"),
  1484 => (x"c1",x"c2",x"55",x"e0"),
  1485 => (x"7d",x"97",x"c0",x"55"),
  1486 => (x"6e",x"49",x"66",x"d4"),
  1487 => (x"87",x"db",x"05",x"a9"),
  1488 => (x"c8",x"48",x"66",x"c4"),
  1489 => (x"ca",x"04",x"a8",x"66"),
  1490 => (x"48",x"66",x"c4",x"87"),
  1491 => (x"a6",x"c8",x"80",x"c1"),
  1492 => (x"c8",x"87",x"c8",x"58"),
  1493 => (x"88",x"c1",x"48",x"66"),
  1494 => (x"e1",x"58",x"a6",x"cc"),
  1495 => (x"4c",x"70",x"87",x"f1"),
  1496 => (x"05",x"ac",x"d0",x"c1"),
  1497 => (x"66",x"d0",x"87",x"c8"),
  1498 => (x"d4",x"80",x"c1",x"48"),
  1499 => (x"d0",x"c1",x"58",x"a6"),
  1500 => (x"e9",x"fd",x"02",x"ac"),
  1501 => (x"a6",x"e0",x"c0",x"87"),
  1502 => (x"78",x"66",x"d4",x"48"),
  1503 => (x"c0",x"48",x"66",x"dc"),
  1504 => (x"05",x"a8",x"66",x"e0"),
  1505 => (x"c0",x"87",x"ca",x"c9"),
  1506 => (x"c0",x"48",x"a6",x"e4"),
  1507 => (x"48",x"74",x"7e",x"78"),
  1508 => (x"c0",x"88",x"fb",x"c0"),
  1509 => (x"70",x"58",x"a6",x"ec"),
  1510 => (x"cf",x"c8",x"02",x"98"),
  1511 => (x"88",x"cb",x"48",x"87"),
  1512 => (x"58",x"a6",x"ec",x"c0"),
  1513 => (x"c1",x"02",x"98",x"70"),
  1514 => (x"c9",x"48",x"87",x"d2"),
  1515 => (x"a6",x"ec",x"c0",x"88"),
  1516 => (x"02",x"98",x"70",x"58"),
  1517 => (x"48",x"87",x"db",x"c3"),
  1518 => (x"ec",x"c0",x"88",x"c4"),
  1519 => (x"98",x"70",x"58",x"a6"),
  1520 => (x"48",x"87",x"d0",x"02"),
  1521 => (x"ec",x"c0",x"88",x"c1"),
  1522 => (x"98",x"70",x"58",x"a6"),
  1523 => (x"87",x"c2",x"c3",x"02"),
  1524 => (x"d8",x"87",x"d3",x"c7"),
  1525 => (x"f0",x"c0",x"48",x"a6"),
  1526 => (x"f2",x"df",x"ff",x"78"),
  1527 => (x"c0",x"4c",x"70",x"87"),
  1528 => (x"c0",x"02",x"ac",x"ec"),
  1529 => (x"a6",x"dc",x"87",x"c3"),
  1530 => (x"ac",x"ec",x"c0",x"5c"),
  1531 => (x"ff",x"87",x"cd",x"02"),
  1532 => (x"70",x"87",x"dc",x"df"),
  1533 => (x"ac",x"ec",x"c0",x"4c"),
  1534 => (x"87",x"f3",x"ff",x"05"),
  1535 => (x"02",x"ac",x"ec",x"c0"),
  1536 => (x"ff",x"87",x"c4",x"c0"),
  1537 => (x"d8",x"87",x"c8",x"df"),
  1538 => (x"66",x"d4",x"1e",x"66"),
  1539 => (x"66",x"d4",x"1e",x"49"),
  1540 => (x"ef",x"c1",x"1e",x"49"),
  1541 => (x"66",x"d4",x"1e",x"c6"),
  1542 => (x"87",x"cb",x"f7",x"49"),
  1543 => (x"1e",x"ca",x"1e",x"c0"),
  1544 => (x"cb",x"49",x"66",x"dc"),
  1545 => (x"66",x"d8",x"c1",x"91"),
  1546 => (x"48",x"a6",x"d8",x"81"),
  1547 => (x"d8",x"78",x"a1",x"c4"),
  1548 => (x"ff",x"49",x"bf",x"66"),
  1549 => (x"d8",x"87",x"dc",x"df"),
  1550 => (x"a8",x"b7",x"c0",x"86"),
  1551 => (x"87",x"c5",x"c1",x"06"),
  1552 => (x"1e",x"de",x"1e",x"c1"),
  1553 => (x"49",x"bf",x"66",x"c8"),
  1554 => (x"87",x"c7",x"df",x"ff"),
  1555 => (x"49",x"70",x"86",x"c8"),
  1556 => (x"88",x"08",x"c0",x"48"),
  1557 => (x"c0",x"58",x"a6",x"dc"),
  1558 => (x"c0",x"06",x"a8",x"b7"),
  1559 => (x"66",x"d8",x"87",x"e7"),
  1560 => (x"a8",x"b7",x"dd",x"48"),
  1561 => (x"6e",x"87",x"de",x"03"),
  1562 => (x"66",x"d8",x"49",x"bf"),
  1563 => (x"51",x"e0",x"c0",x"81"),
  1564 => (x"c1",x"49",x"66",x"d8"),
  1565 => (x"81",x"bf",x"6e",x"81"),
  1566 => (x"d8",x"51",x"c1",x"c2"),
  1567 => (x"81",x"c2",x"49",x"66"),
  1568 => (x"c0",x"81",x"bf",x"6e"),
  1569 => (x"48",x"66",x"cc",x"51"),
  1570 => (x"a6",x"d0",x"80",x"c1"),
  1571 => (x"c4",x"7e",x"c1",x"58"),
  1572 => (x"df",x"ff",x"87",x"da"),
  1573 => (x"a6",x"dc",x"87",x"ec"),
  1574 => (x"e5",x"df",x"ff",x"58"),
  1575 => (x"a6",x"ec",x"c0",x"87"),
  1576 => (x"a8",x"ec",x"c0",x"58"),
  1577 => (x"87",x"ca",x"c0",x"05"),
  1578 => (x"48",x"a6",x"e8",x"c0"),
  1579 => (x"c0",x"78",x"66",x"d8"),
  1580 => (x"dc",x"ff",x"87",x"c4"),
  1581 => (x"66",x"c4",x"87",x"d9"),
  1582 => (x"c1",x"91",x"cb",x"49"),
  1583 => (x"71",x"48",x"66",x"c0"),
  1584 => (x"6e",x"7e",x"70",x"80"),
  1585 => (x"6e",x"82",x"c8",x"4a"),
  1586 => (x"d8",x"81",x"ca",x"49"),
  1587 => (x"e8",x"c0",x"51",x"66"),
  1588 => (x"81",x"c1",x"49",x"66"),
  1589 => (x"c1",x"89",x"66",x"d8"),
  1590 => (x"70",x"30",x"71",x"48"),
  1591 => (x"71",x"89",x"c1",x"49"),
  1592 => (x"ca",x"c4",x"7a",x"97"),
  1593 => (x"d8",x"49",x"bf",x"e1"),
  1594 => (x"6a",x"97",x"29",x"66"),
  1595 => (x"98",x"71",x"48",x"4a"),
  1596 => (x"58",x"a6",x"f0",x"c0"),
  1597 => (x"81",x"c4",x"49",x"6e"),
  1598 => (x"e0",x"c0",x"4d",x"69"),
  1599 => (x"66",x"dc",x"48",x"66"),
  1600 => (x"c8",x"c0",x"02",x"a8"),
  1601 => (x"48",x"a6",x"d8",x"87"),
  1602 => (x"c5",x"c0",x"78",x"c0"),
  1603 => (x"48",x"a6",x"d8",x"87"),
  1604 => (x"66",x"d8",x"78",x"c1"),
  1605 => (x"1e",x"e0",x"c0",x"1e"),
  1606 => (x"db",x"ff",x"49",x"75"),
  1607 => (x"86",x"c8",x"87",x"f5"),
  1608 => (x"b7",x"c0",x"4c",x"70"),
  1609 => (x"d4",x"c1",x"06",x"ac"),
  1610 => (x"c0",x"85",x"74",x"87"),
  1611 => (x"89",x"74",x"49",x"e0"),
  1612 => (x"e8",x"c1",x"4b",x"75"),
  1613 => (x"fe",x"71",x"4a",x"f8"),
  1614 => (x"c2",x"87",x"fe",x"dd"),
  1615 => (x"66",x"e4",x"c0",x"85"),
  1616 => (x"c0",x"80",x"c1",x"48"),
  1617 => (x"c0",x"58",x"a6",x"e8"),
  1618 => (x"c1",x"49",x"66",x"ec"),
  1619 => (x"02",x"a9",x"70",x"81"),
  1620 => (x"d8",x"87",x"c8",x"c0"),
  1621 => (x"78",x"c0",x"48",x"a6"),
  1622 => (x"d8",x"87",x"c5",x"c0"),
  1623 => (x"78",x"c1",x"48",x"a6"),
  1624 => (x"c2",x"1e",x"66",x"d8"),
  1625 => (x"e0",x"c0",x"49",x"a4"),
  1626 => (x"70",x"88",x"71",x"48"),
  1627 => (x"49",x"75",x"1e",x"49"),
  1628 => (x"87",x"df",x"da",x"ff"),
  1629 => (x"b7",x"c0",x"86",x"c8"),
  1630 => (x"c0",x"ff",x"01",x"a8"),
  1631 => (x"66",x"e4",x"c0",x"87"),
  1632 => (x"87",x"d1",x"c0",x"02"),
  1633 => (x"81",x"c9",x"49",x"6e"),
  1634 => (x"51",x"66",x"e4",x"c0"),
  1635 => (x"d4",x"c1",x"48",x"6e"),
  1636 => (x"cc",x"c0",x"78",x"d3"),
  1637 => (x"c9",x"49",x"6e",x"87"),
  1638 => (x"6e",x"51",x"c2",x"81"),
  1639 => (x"c7",x"d5",x"c1",x"48"),
  1640 => (x"c0",x"7e",x"c1",x"78"),
  1641 => (x"d9",x"ff",x"87",x"c6"),
  1642 => (x"4c",x"70",x"87",x"d5"),
  1643 => (x"f5",x"c0",x"02",x"6e"),
  1644 => (x"48",x"66",x"c4",x"87"),
  1645 => (x"04",x"a8",x"66",x"c8"),
  1646 => (x"c4",x"87",x"cb",x"c0"),
  1647 => (x"80",x"c1",x"48",x"66"),
  1648 => (x"c0",x"58",x"a6",x"c8"),
  1649 => (x"66",x"c8",x"87",x"e0"),
  1650 => (x"cc",x"88",x"c1",x"48"),
  1651 => (x"d5",x"c0",x"58",x"a6"),
  1652 => (x"ac",x"c6",x"c1",x"87"),
  1653 => (x"87",x"c8",x"c0",x"05"),
  1654 => (x"c1",x"48",x"66",x"cc"),
  1655 => (x"58",x"a6",x"d0",x"80"),
  1656 => (x"87",x"db",x"d8",x"ff"),
  1657 => (x"66",x"d0",x"4c",x"70"),
  1658 => (x"d4",x"80",x"c1",x"48"),
  1659 => (x"9c",x"74",x"58",x"a6"),
  1660 => (x"87",x"cb",x"c0",x"02"),
  1661 => (x"c1",x"48",x"66",x"c4"),
  1662 => (x"04",x"a8",x"66",x"c8"),
  1663 => (x"ff",x"87",x"ca",x"f3"),
  1664 => (x"c4",x"87",x"f3",x"d7"),
  1665 => (x"a8",x"c7",x"48",x"66"),
  1666 => (x"87",x"e5",x"c0",x"03"),
  1667 => (x"48",x"f4",x"c6",x"c4"),
  1668 => (x"66",x"c4",x"78",x"c0"),
  1669 => (x"c1",x"91",x"cb",x"49"),
  1670 => (x"c4",x"81",x"66",x"c0"),
  1671 => (x"4a",x"6a",x"4a",x"a1"),
  1672 => (x"c4",x"79",x"52",x"c0"),
  1673 => (x"80",x"c1",x"48",x"66"),
  1674 => (x"c7",x"58",x"a6",x"c8"),
  1675 => (x"db",x"ff",x"04",x"a8"),
  1676 => (x"8e",x"d0",x"ff",x"87"),
  1677 => (x"87",x"d9",x"de",x"ff"),
  1678 => (x"1e",x"00",x"20",x"3a"),
  1679 => (x"4b",x"71",x"1e",x"73"),
  1680 => (x"87",x"c6",x"02",x"9b"),
  1681 => (x"48",x"f0",x"c6",x"c4"),
  1682 => (x"1e",x"c7",x"78",x"c0"),
  1683 => (x"bf",x"f0",x"c6",x"c4"),
  1684 => (x"ed",x"c1",x"1e",x"49"),
  1685 => (x"c6",x"c4",x"1e",x"d3"),
  1686 => (x"ee",x"49",x"bf",x"ec"),
  1687 => (x"86",x"cc",x"87",x"fe"),
  1688 => (x"bf",x"ec",x"c6",x"c4"),
  1689 => (x"87",x"c3",x"ea",x"49"),
  1690 => (x"c8",x"02",x"9b",x"73"),
  1691 => (x"d3",x"ed",x"c1",x"87"),
  1692 => (x"db",x"e7",x"c0",x"49"),
  1693 => (x"dc",x"dd",x"ff",x"87"),
  1694 => (x"1e",x"73",x"1e",x"87"),
  1695 => (x"f7",x"c3",x"4b",x"c0"),
  1696 => (x"50",x"c0",x"48",x"eb"),
  1697 => (x"bf",x"f6",x"ee",x"c1"),
  1698 => (x"e6",x"c8",x"c2",x"49"),
  1699 => (x"05",x"98",x"70",x"87"),
  1700 => (x"ea",x"c1",x"87",x"c4"),
  1701 => (x"48",x"73",x"4b",x"dc"),
  1702 => (x"87",x"f9",x"dc",x"ff"),
  1703 => (x"20",x"4d",x"4f",x"52"),
  1704 => (x"64",x"61",x"6f",x"6c"),
  1705 => (x"20",x"67",x"6e",x"69"),
  1706 => (x"6c",x"69",x"61",x"66"),
  1707 => (x"1e",x"00",x"64",x"65"),
  1708 => (x"c1",x"87",x"f2",x"c7"),
  1709 => (x"87",x"c3",x"fe",x"49"),
  1710 => (x"87",x"fe",x"e6",x"fe"),
  1711 => (x"cd",x"02",x"98",x"70"),
  1712 => (x"fb",x"ef",x"fe",x"87"),
  1713 => (x"02",x"98",x"70",x"87"),
  1714 => (x"4a",x"c1",x"87",x"c4"),
  1715 => (x"4a",x"c0",x"87",x"c2"),
  1716 => (x"ce",x"05",x"9a",x"72"),
  1717 => (x"c1",x"1e",x"c0",x"87"),
  1718 => (x"c0",x"49",x"c3",x"ec"),
  1719 => (x"c4",x"87",x"c1",x"f3"),
  1720 => (x"c2",x"87",x"fe",x"86"),
  1721 => (x"c0",x"87",x"ee",x"cc"),
  1722 => (x"ce",x"ec",x"c1",x"1e"),
  1723 => (x"ef",x"f2",x"c0",x"49"),
  1724 => (x"fe",x"1e",x"c0",x"87"),
  1725 => (x"49",x"70",x"87",x"c3"),
  1726 => (x"87",x"e4",x"f2",x"c0"),
  1727 => (x"f8",x"87",x"e5",x"c3"),
  1728 => (x"53",x"4f",x"26",x"8e"),
  1729 => (x"61",x"66",x"20",x"44"),
  1730 => (x"64",x"65",x"6c",x"69"),
  1731 => (x"6f",x"42",x"00",x"2e"),
  1732 => (x"6e",x"69",x"74",x"6f"),
  1733 => (x"2e",x"2e",x"2e",x"67"),
  1734 => (x"fc",x"c1",x"1e",x"00"),
  1735 => (x"e9",x"c0",x"87",x"c2"),
  1736 => (x"fb",x"c1",x"87",x"cc"),
  1737 => (x"c0",x"c2",x"87",x"fa"),
  1738 => (x"87",x"ee",x"87",x"f8"),
  1739 => (x"c4",x"1e",x"4f",x"26"),
  1740 => (x"c0",x"48",x"f0",x"c6"),
  1741 => (x"ec",x"c6",x"c4",x"78"),
  1742 => (x"fd",x"78",x"c0",x"48"),
  1743 => (x"d8",x"ff",x"87",x"f1"),
  1744 => (x"26",x"48",x"c0",x"87"),
  1745 => (x"45",x"20",x"80",x"4f"),
  1746 => (x"00",x"74",x"69",x"78"),
  1747 => (x"61",x"42",x"20",x"80"),
  1748 => (x"c3",x"00",x"6b",x"63"),
  1749 => (x"c5",x"00",x"00",x"14"),
  1750 => (x"00",x"00",x"00",x"41"),
  1751 => (x"14",x"c3",x"00",x"00"),
  1752 => (x"41",x"e3",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"14",x"c3",x"00"),
  1755 => (x"00",x"42",x"01",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"14",x"c3"),
  1758 => (x"00",x"00",x"42",x"1f"),
  1759 => (x"c3",x"00",x"00",x"00"),
  1760 => (x"3d",x"00",x"00",x"14"),
  1761 => (x"00",x"00",x"00",x"42"),
  1762 => (x"14",x"c3",x"00",x"00"),
  1763 => (x"42",x"5b",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"14",x"c3",x"00"),
  1766 => (x"00",x"42",x"79",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"14",x"c3"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"58",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"15"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"1b",x"ba",x"00",x"00"),
  1774 => (x"45",x"4e",x"00",x"00"),
  1775 => (x"4f",x"45",x"47",x"4f"),
  1776 => (x"4f",x"52",x"20",x"20"),
  1777 => (x"6f",x"4c",x"00",x"4d"),
  1778 => (x"2a",x"20",x"64",x"61"),
  1779 => (x"fe",x"1e",x"00",x"2e"),
  1780 => (x"78",x"c0",x"48",x"f0"),
  1781 => (x"09",x"79",x"09",x"cd"),
  1782 => (x"1e",x"1e",x"4f",x"26"),
  1783 => (x"7e",x"bf",x"f0",x"fe"),
  1784 => (x"4f",x"26",x"26",x"48"),
  1785 => (x"48",x"f0",x"fe",x"1e"),
  1786 => (x"4f",x"26",x"78",x"c1"),
  1787 => (x"48",x"f0",x"fe",x"1e"),
  1788 => (x"4f",x"26",x"78",x"c0"),
  1789 => (x"c0",x"4a",x"71",x"1e"),
  1790 => (x"4f",x"26",x"52",x"52"),
  1791 => (x"5c",x"5b",x"5e",x"0e"),
  1792 => (x"86",x"f4",x"0e",x"5d"),
  1793 => (x"6d",x"97",x"4d",x"71"),
  1794 => (x"4c",x"a5",x"c1",x"7e"),
  1795 => (x"c8",x"48",x"6c",x"97"),
  1796 => (x"48",x"6e",x"58",x"a6"),
  1797 => (x"05",x"a8",x"66",x"c4"),
  1798 => (x"48",x"ff",x"87",x"c5"),
  1799 => (x"ff",x"87",x"e6",x"c0"),
  1800 => (x"a5",x"c2",x"87",x"ca"),
  1801 => (x"4b",x"6c",x"97",x"49"),
  1802 => (x"97",x"4b",x"a3",x"71"),
  1803 => (x"6c",x"97",x"4b",x"6b"),
  1804 => (x"c1",x"48",x"6e",x"7e"),
  1805 => (x"58",x"a6",x"c8",x"80"),
  1806 => (x"a6",x"cc",x"98",x"c7"),
  1807 => (x"7c",x"97",x"70",x"58"),
  1808 => (x"73",x"87",x"e1",x"fe"),
  1809 => (x"26",x"8e",x"f4",x"48"),
  1810 => (x"26",x"4c",x"26",x"4d"),
  1811 => (x"0e",x"4f",x"26",x"4b"),
  1812 => (x"0e",x"5c",x"5b",x"5e"),
  1813 => (x"4c",x"71",x"86",x"f4"),
  1814 => (x"c3",x"4a",x"66",x"d8"),
  1815 => (x"a4",x"c2",x"9a",x"ff"),
  1816 => (x"49",x"6c",x"97",x"4b"),
  1817 => (x"72",x"49",x"a1",x"73"),
  1818 => (x"7e",x"6c",x"97",x"51"),
  1819 => (x"80",x"c1",x"48",x"6e"),
  1820 => (x"c7",x"58",x"a6",x"c8"),
  1821 => (x"58",x"a6",x"cc",x"98"),
  1822 => (x"8e",x"f4",x"54",x"70"),
  1823 => (x"1e",x"87",x"ca",x"ff"),
  1824 => (x"87",x"e8",x"fd",x"1e"),
  1825 => (x"49",x"4a",x"bf",x"e0"),
  1826 => (x"99",x"c0",x"e0",x"c0"),
  1827 => (x"72",x"87",x"cb",x"02"),
  1828 => (x"d7",x"ca",x"c4",x"1e"),
  1829 => (x"87",x"f7",x"fe",x"49"),
  1830 => (x"fd",x"fc",x"86",x"c4"),
  1831 => (x"fd",x"7e",x"70",x"87"),
  1832 => (x"26",x"26",x"87",x"c2"),
  1833 => (x"ca",x"c4",x"1e",x"4f"),
  1834 => (x"c7",x"fd",x"49",x"d7"),
  1835 => (x"ff",x"f1",x"c1",x"87"),
  1836 => (x"87",x"da",x"fc",x"49"),
  1837 => (x"26",x"87",x"d5",x"c6"),
  1838 => (x"5b",x"5e",x"0e",x"4f"),
  1839 => (x"c4",x"0e",x"5d",x"5c"),
  1840 => (x"4a",x"bf",x"f6",x"ca"),
  1841 => (x"bf",x"cd",x"f4",x"c1"),
  1842 => (x"bc",x"72",x"4c",x"49"),
  1843 => (x"db",x"fc",x"4d",x"71"),
  1844 => (x"74",x"4b",x"c0",x"87"),
  1845 => (x"02",x"99",x"d0",x"49"),
  1846 => (x"49",x"75",x"87",x"d5"),
  1847 => (x"1e",x"71",x"99",x"d0"),
  1848 => (x"fb",x"c1",x"1e",x"c0"),
  1849 => (x"82",x"73",x"4a",x"db"),
  1850 => (x"ca",x"c1",x"49",x"12"),
  1851 => (x"c1",x"86",x"c8",x"87"),
  1852 => (x"c8",x"83",x"2d",x"2c"),
  1853 => (x"da",x"ff",x"04",x"ab"),
  1854 => (x"87",x"e8",x"fb",x"87"),
  1855 => (x"48",x"cd",x"f4",x"c1"),
  1856 => (x"bf",x"f6",x"ca",x"c4"),
  1857 => (x"26",x"4d",x"26",x"78"),
  1858 => (x"26",x"4b",x"26",x"4c"),
  1859 => (x"00",x"00",x"00",x"4f"),
  1860 => (x"1e",x"73",x"1e",x"00"),
  1861 => (x"4a",x"c0",x"4b",x"71"),
  1862 => (x"49",x"db",x"fb",x"c1"),
  1863 => (x"69",x"97",x"81",x"72"),
  1864 => (x"05",x"a9",x"73",x"49"),
  1865 => (x"48",x"c1",x"87",x"c4"),
  1866 => (x"82",x"c1",x"87",x"ca"),
  1867 => (x"04",x"aa",x"b7",x"c8"),
  1868 => (x"48",x"c0",x"87",x"e6"),
  1869 => (x"1e",x"87",x"d2",x"ff"),
  1870 => (x"4b",x"71",x"1e",x"73"),
  1871 => (x"87",x"d1",x"ff",x"49"),
  1872 => (x"c0",x"02",x"98",x"70"),
  1873 => (x"d0",x"ff",x"87",x"ec"),
  1874 => (x"78",x"e1",x"c8",x"48"),
  1875 => (x"c5",x"48",x"d4",x"ff"),
  1876 => (x"02",x"66",x"c8",x"78"),
  1877 => (x"e0",x"c3",x"87",x"c3"),
  1878 => (x"02",x"66",x"cc",x"78"),
  1879 => (x"d4",x"ff",x"87",x"c6"),
  1880 => (x"78",x"f0",x"c3",x"48"),
  1881 => (x"73",x"48",x"d4",x"ff"),
  1882 => (x"48",x"d0",x"ff",x"78"),
  1883 => (x"c0",x"78",x"e1",x"c8"),
  1884 => (x"d4",x"fe",x"78",x"e0"),
  1885 => (x"5b",x"5e",x"0e",x"87"),
  1886 => (x"4c",x"71",x"0e",x"5c"),
  1887 => (x"49",x"d7",x"ca",x"c4"),
  1888 => (x"70",x"87",x"f9",x"f9"),
  1889 => (x"aa",x"b7",x"c0",x"4a"),
  1890 => (x"87",x"e3",x"c2",x"04"),
  1891 => (x"05",x"aa",x"e0",x"c3"),
  1892 => (x"f8",x"c1",x"87",x"c9"),
  1893 => (x"78",x"c1",x"48",x"f8"),
  1894 => (x"c3",x"87",x"d4",x"c2"),
  1895 => (x"c9",x"05",x"aa",x"f0"),
  1896 => (x"f4",x"f8",x"c1",x"87"),
  1897 => (x"c1",x"78",x"c1",x"48"),
  1898 => (x"f8",x"c1",x"87",x"f5"),
  1899 => (x"c7",x"02",x"bf",x"f8"),
  1900 => (x"c2",x"4b",x"72",x"87"),
  1901 => (x"87",x"c2",x"b3",x"c0"),
  1902 => (x"9c",x"74",x"4b",x"72"),
  1903 => (x"c1",x"87",x"d1",x"05"),
  1904 => (x"1e",x"bf",x"f4",x"f8"),
  1905 => (x"bf",x"f8",x"f8",x"c1"),
  1906 => (x"fd",x"49",x"72",x"1e"),
  1907 => (x"86",x"c8",x"87",x"e9"),
  1908 => (x"bf",x"f4",x"f8",x"c1"),
  1909 => (x"87",x"e0",x"c0",x"02"),
  1910 => (x"b7",x"c4",x"49",x"73"),
  1911 => (x"fa",x"c1",x"91",x"29"),
  1912 => (x"4a",x"73",x"81",x"db"),
  1913 => (x"92",x"c2",x"9a",x"cf"),
  1914 => (x"30",x"72",x"48",x"c1"),
  1915 => (x"ba",x"ff",x"4a",x"70"),
  1916 => (x"98",x"69",x"48",x"72"),
  1917 => (x"87",x"db",x"79",x"70"),
  1918 => (x"b7",x"c4",x"49",x"73"),
  1919 => (x"fa",x"c1",x"91",x"29"),
  1920 => (x"4a",x"73",x"81",x"db"),
  1921 => (x"92",x"c2",x"9a",x"cf"),
  1922 => (x"30",x"72",x"48",x"c3"),
  1923 => (x"69",x"48",x"4a",x"70"),
  1924 => (x"c1",x"79",x"70",x"b0"),
  1925 => (x"c0",x"48",x"f8",x"f8"),
  1926 => (x"f4",x"f8",x"c1",x"78"),
  1927 => (x"c4",x"78",x"c0",x"48"),
  1928 => (x"f7",x"49",x"d7",x"ca"),
  1929 => (x"4a",x"70",x"87",x"d6"),
  1930 => (x"03",x"aa",x"b7",x"c0"),
  1931 => (x"c0",x"87",x"dd",x"fd"),
  1932 => (x"87",x"d3",x"fb",x"48"),
  1933 => (x"00",x"00",x"00",x"00"),
  1934 => (x"00",x"00",x"00",x"00"),
  1935 => (x"71",x"1e",x"73",x"1e"),
  1936 => (x"87",x"f5",x"f9",x"4b"),
  1937 => (x"ec",x"fc",x"49",x"73"),
  1938 => (x"87",x"fd",x"fa",x"87"),
  1939 => (x"72",x"4a",x"c0",x"1e"),
  1940 => (x"c1",x"91",x"c4",x"49"),
  1941 => (x"c0",x"81",x"db",x"fa"),
  1942 => (x"d0",x"82",x"c1",x"79"),
  1943 => (x"ee",x"04",x"aa",x"b7"),
  1944 => (x"0e",x"4f",x"26",x"87"),
  1945 => (x"5d",x"5c",x"5b",x"5e"),
  1946 => (x"f5",x"4d",x"71",x"0e"),
  1947 => (x"4a",x"75",x"87",x"fe"),
  1948 => (x"92",x"2a",x"b7",x"c4"),
  1949 => (x"82",x"db",x"fa",x"c1"),
  1950 => (x"9c",x"cf",x"4c",x"75"),
  1951 => (x"49",x"6a",x"94",x"c2"),
  1952 => (x"c3",x"2b",x"74",x"4b"),
  1953 => (x"74",x"48",x"c2",x"9b"),
  1954 => (x"ff",x"4c",x"70",x"30"),
  1955 => (x"71",x"48",x"74",x"bc"),
  1956 => (x"f5",x"7a",x"70",x"98"),
  1957 => (x"48",x"73",x"87",x"ce"),
  1958 => (x"00",x"87",x"ea",x"f9"),
  1959 => (x"00",x"00",x"00",x"00"),
  1960 => (x"00",x"00",x"00",x"00"),
  1961 => (x"00",x"00",x"00",x"00"),
  1962 => (x"00",x"00",x"00",x"00"),
  1963 => (x"00",x"00",x"00",x"00"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"00",x"00"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"00"),
  1969 => (x"00",x"00",x"00",x"00"),
  1970 => (x"00",x"00",x"00",x"00"),
  1971 => (x"00",x"00",x"00",x"00"),
  1972 => (x"00",x"00",x"00",x"00"),
  1973 => (x"00",x"00",x"00",x"00"),
  1974 => (x"16",x"00",x"00",x"00"),
  1975 => (x"2e",x"25",x"26",x"1e"),
  1976 => (x"1e",x"3e",x"3d",x"36"),
  1977 => (x"c8",x"48",x"d0",x"ff"),
  1978 => (x"48",x"71",x"78",x"e1"),
  1979 => (x"78",x"08",x"d4",x"ff"),
  1980 => (x"ff",x"1e",x"4f",x"26"),
  1981 => (x"e1",x"c8",x"48",x"d0"),
  1982 => (x"ff",x"48",x"71",x"78"),
  1983 => (x"c4",x"78",x"08",x"d4"),
  1984 => (x"d4",x"ff",x"48",x"66"),
  1985 => (x"4f",x"26",x"78",x"08"),
  1986 => (x"c4",x"4a",x"71",x"1e"),
  1987 => (x"72",x"1e",x"49",x"66"),
  1988 => (x"87",x"de",x"ff",x"49"),
  1989 => (x"c0",x"48",x"d0",x"ff"),
  1990 => (x"26",x"26",x"78",x"e0"),
  1991 => (x"4a",x"71",x"1e",x"4f"),
  1992 => (x"c1",x"1e",x"66",x"c4"),
  1993 => (x"ff",x"49",x"a2",x"e0"),
  1994 => (x"66",x"c8",x"87",x"c8"),
  1995 => (x"29",x"b7",x"c8",x"49"),
  1996 => (x"71",x"48",x"d4",x"ff"),
  1997 => (x"48",x"d0",x"ff",x"78"),
  1998 => (x"26",x"78",x"e0",x"c0"),
  1999 => (x"ff",x"1e",x"4f",x"26"),
  2000 => (x"ff",x"c3",x"4a",x"d4"),
  2001 => (x"48",x"d0",x"ff",x"7a"),
  2002 => (x"de",x"78",x"e1",x"c8"),
  2003 => (x"e1",x"ca",x"c4",x"7a"),
  2004 => (x"48",x"49",x"7a",x"bf"),
  2005 => (x"7a",x"70",x"28",x"c8"),
  2006 => (x"28",x"d0",x"48",x"71"),
  2007 => (x"48",x"71",x"7a",x"70"),
  2008 => (x"7a",x"70",x"28",x"d8"),
  2009 => (x"c0",x"48",x"d0",x"ff"),
  2010 => (x"4f",x"26",x"78",x"e0"),
  2011 => (x"5c",x"5b",x"5e",x"0e"),
  2012 => (x"4c",x"71",x"0e",x"5d"),
  2013 => (x"bf",x"e1",x"ca",x"c4"),
  2014 => (x"2b",x"74",x"4b",x"4d"),
  2015 => (x"c1",x"9b",x"66",x"d0"),
  2016 => (x"ab",x"66",x"d4",x"83"),
  2017 => (x"c0",x"87",x"c2",x"04"),
  2018 => (x"d0",x"4a",x"74",x"4b"),
  2019 => (x"31",x"72",x"49",x"66"),
  2020 => (x"99",x"75",x"b9",x"ff"),
  2021 => (x"30",x"72",x"48",x"73"),
  2022 => (x"71",x"48",x"4a",x"70"),
  2023 => (x"e5",x"ca",x"c4",x"b0"),
  2024 => (x"87",x"da",x"fe",x"58"),
  2025 => (x"4c",x"26",x"4d",x"26"),
  2026 => (x"4f",x"26",x"4b",x"26"),
  2027 => (x"48",x"d0",x"ff",x"1e"),
  2028 => (x"71",x"78",x"c9",x"c8"),
  2029 => (x"08",x"d4",x"ff",x"48"),
  2030 => (x"1e",x"4f",x"26",x"78"),
  2031 => (x"eb",x"49",x"4a",x"71"),
  2032 => (x"48",x"d0",x"ff",x"87"),
  2033 => (x"4f",x"26",x"78",x"c8"),
  2034 => (x"71",x"1e",x"73",x"1e"),
  2035 => (x"f1",x"ca",x"c4",x"4b"),
  2036 => (x"87",x"c3",x"02",x"bf"),
  2037 => (x"ff",x"87",x"eb",x"c2"),
  2038 => (x"c9",x"c8",x"48",x"d0"),
  2039 => (x"c0",x"49",x"73",x"78"),
  2040 => (x"d4",x"ff",x"b1",x"e0"),
  2041 => (x"c4",x"78",x"71",x"48"),
  2042 => (x"c0",x"48",x"e5",x"ca"),
  2043 => (x"02",x"66",x"c8",x"78"),
  2044 => (x"ff",x"c3",x"87",x"c5"),
  2045 => (x"c0",x"87",x"c2",x"49"),
  2046 => (x"ed",x"ca",x"c4",x"49"),
  2047 => (x"02",x"66",x"cc",x"59"),
  2048 => (x"d5",x"c5",x"87",x"c6"),
  2049 => (x"87",x"c4",x"4a",x"d5"),
  2050 => (x"4a",x"ff",x"ff",x"cf"),
  2051 => (x"5a",x"f1",x"ca",x"c4"),
  2052 => (x"48",x"f1",x"ca",x"c4"),
  2053 => (x"87",x"c4",x"78",x"c1"),
  2054 => (x"4c",x"26",x"4d",x"26"),
  2055 => (x"4f",x"26",x"4b",x"26"),
  2056 => (x"5c",x"5b",x"5e",x"0e"),
  2057 => (x"4a",x"71",x"0e",x"5d"),
  2058 => (x"bf",x"ed",x"ca",x"c4"),
  2059 => (x"02",x"9a",x"72",x"4c"),
  2060 => (x"c8",x"49",x"87",x"cb"),
  2061 => (x"fe",x"fe",x"c1",x"91"),
  2062 => (x"c4",x"83",x"71",x"4b"),
  2063 => (x"fe",x"c2",x"c2",x"87"),
  2064 => (x"13",x"4d",x"c0",x"4b"),
  2065 => (x"c4",x"99",x"74",x"49"),
  2066 => (x"b9",x"bf",x"e9",x"ca"),
  2067 => (x"71",x"48",x"d4",x"ff"),
  2068 => (x"2c",x"b7",x"c1",x"78"),
  2069 => (x"ad",x"b7",x"c8",x"85"),
  2070 => (x"c4",x"87",x"e8",x"04"),
  2071 => (x"48",x"bf",x"e5",x"ca"),
  2072 => (x"ca",x"c4",x"80",x"c8"),
  2073 => (x"ef",x"fe",x"58",x"e9"),
  2074 => (x"1e",x"73",x"1e",x"87"),
  2075 => (x"4a",x"13",x"4b",x"71"),
  2076 => (x"87",x"cb",x"02",x"9a"),
  2077 => (x"e7",x"fe",x"49",x"72"),
  2078 => (x"9a",x"4a",x"13",x"87"),
  2079 => (x"fe",x"87",x"f5",x"05"),
  2080 => (x"c4",x"1e",x"87",x"da"),
  2081 => (x"49",x"bf",x"e5",x"ca"),
  2082 => (x"48",x"e5",x"ca",x"c4"),
  2083 => (x"c4",x"78",x"a1",x"c1"),
  2084 => (x"03",x"a9",x"b7",x"c0"),
  2085 => (x"d4",x"ff",x"87",x"db"),
  2086 => (x"e9",x"ca",x"c4",x"48"),
  2087 => (x"ca",x"c4",x"78",x"bf"),
  2088 => (x"c4",x"49",x"bf",x"e5"),
  2089 => (x"c1",x"48",x"e5",x"ca"),
  2090 => (x"c0",x"c4",x"78",x"a1"),
  2091 => (x"e5",x"04",x"a9",x"b7"),
  2092 => (x"48",x"d0",x"ff",x"87"),
  2093 => (x"ca",x"c4",x"78",x"c8"),
  2094 => (x"78",x"c0",x"48",x"f1"),
  2095 => (x"00",x"00",x"4f",x"26"),
  2096 => (x"00",x"00",x"00",x"00"),
  2097 => (x"00",x"00",x"00",x"00"),
  2098 => (x"00",x"5f",x"5f",x"00"),
  2099 => (x"03",x"00",x"00",x"00"),
  2100 => (x"03",x"03",x"00",x"03"),
  2101 => (x"7f",x"14",x"00",x"00"),
  2102 => (x"7f",x"7f",x"14",x"7f"),
  2103 => (x"24",x"00",x"00",x"14"),
  2104 => (x"3a",x"6b",x"6b",x"2e"),
  2105 => (x"6a",x"4c",x"00",x"12"),
  2106 => (x"56",x"6c",x"18",x"36"),
  2107 => (x"7e",x"30",x"00",x"32"),
  2108 => (x"3a",x"77",x"59",x"4f"),
  2109 => (x"00",x"00",x"40",x"68"),
  2110 => (x"00",x"03",x"07",x"04"),
  2111 => (x"00",x"00",x"00",x"00"),
  2112 => (x"41",x"63",x"3e",x"1c"),
  2113 => (x"00",x"00",x"00",x"00"),
  2114 => (x"1c",x"3e",x"63",x"41"),
  2115 => (x"2a",x"08",x"00",x"00"),
  2116 => (x"3e",x"1c",x"1c",x"3e"),
  2117 => (x"08",x"00",x"08",x"2a"),
  2118 => (x"08",x"3e",x"3e",x"08"),
  2119 => (x"00",x"00",x"00",x"08"),
  2120 => (x"00",x"60",x"e0",x"80"),
  2121 => (x"08",x"00",x"00",x"00"),
  2122 => (x"08",x"08",x"08",x"08"),
  2123 => (x"00",x"00",x"00",x"08"),
  2124 => (x"00",x"60",x"60",x"00"),
  2125 => (x"60",x"40",x"00",x"00"),
  2126 => (x"06",x"0c",x"18",x"30"),
  2127 => (x"3e",x"00",x"01",x"03"),
  2128 => (x"7f",x"4d",x"59",x"7f"),
  2129 => (x"04",x"00",x"00",x"3e"),
  2130 => (x"00",x"7f",x"7f",x"06"),
  2131 => (x"42",x"00",x"00",x"00"),
  2132 => (x"4f",x"59",x"71",x"63"),
  2133 => (x"22",x"00",x"00",x"46"),
  2134 => (x"7f",x"49",x"49",x"63"),
  2135 => (x"1c",x"18",x"00",x"36"),
  2136 => (x"7f",x"7f",x"13",x"16"),
  2137 => (x"27",x"00",x"00",x"10"),
  2138 => (x"7d",x"45",x"45",x"67"),
  2139 => (x"3c",x"00",x"00",x"39"),
  2140 => (x"79",x"49",x"4b",x"7e"),
  2141 => (x"01",x"00",x"00",x"30"),
  2142 => (x"0f",x"79",x"71",x"01"),
  2143 => (x"36",x"00",x"00",x"07"),
  2144 => (x"7f",x"49",x"49",x"7f"),
  2145 => (x"06",x"00",x"00",x"36"),
  2146 => (x"3f",x"69",x"49",x"4f"),
  2147 => (x"00",x"00",x"00",x"1e"),
  2148 => (x"00",x"66",x"66",x"00"),
  2149 => (x"00",x"00",x"00",x"00"),
  2150 => (x"00",x"66",x"e6",x"80"),
  2151 => (x"08",x"00",x"00",x"00"),
  2152 => (x"22",x"14",x"14",x"08"),
  2153 => (x"14",x"00",x"00",x"22"),
  2154 => (x"14",x"14",x"14",x"14"),
  2155 => (x"22",x"00",x"00",x"14"),
  2156 => (x"08",x"14",x"14",x"22"),
  2157 => (x"02",x"00",x"00",x"08"),
  2158 => (x"0f",x"59",x"51",x"03"),
  2159 => (x"7f",x"3e",x"00",x"06"),
  2160 => (x"1f",x"55",x"5d",x"41"),
  2161 => (x"7e",x"00",x"00",x"1e"),
  2162 => (x"7f",x"09",x"09",x"7f"),
  2163 => (x"7f",x"00",x"00",x"7e"),
  2164 => (x"7f",x"49",x"49",x"7f"),
  2165 => (x"1c",x"00",x"00",x"36"),
  2166 => (x"41",x"41",x"63",x"3e"),
  2167 => (x"7f",x"00",x"00",x"41"),
  2168 => (x"3e",x"63",x"41",x"7f"),
  2169 => (x"7f",x"00",x"00",x"1c"),
  2170 => (x"41",x"49",x"49",x"7f"),
  2171 => (x"7f",x"00",x"00",x"41"),
  2172 => (x"01",x"09",x"09",x"7f"),
  2173 => (x"3e",x"00",x"00",x"01"),
  2174 => (x"7b",x"49",x"41",x"7f"),
  2175 => (x"7f",x"00",x"00",x"7a"),
  2176 => (x"7f",x"08",x"08",x"7f"),
  2177 => (x"00",x"00",x"00",x"7f"),
  2178 => (x"41",x"7f",x"7f",x"41"),
  2179 => (x"20",x"00",x"00",x"00"),
  2180 => (x"7f",x"40",x"40",x"60"),
  2181 => (x"7f",x"7f",x"00",x"3f"),
  2182 => (x"63",x"36",x"1c",x"08"),
  2183 => (x"7f",x"00",x"00",x"41"),
  2184 => (x"40",x"40",x"40",x"7f"),
  2185 => (x"7f",x"7f",x"00",x"40"),
  2186 => (x"7f",x"06",x"0c",x"06"),
  2187 => (x"7f",x"7f",x"00",x"7f"),
  2188 => (x"7f",x"18",x"0c",x"06"),
  2189 => (x"3e",x"00",x"00",x"7f"),
  2190 => (x"7f",x"41",x"41",x"7f"),
  2191 => (x"7f",x"00",x"00",x"3e"),
  2192 => (x"0f",x"09",x"09",x"7f"),
  2193 => (x"7f",x"3e",x"00",x"06"),
  2194 => (x"7e",x"7f",x"61",x"41"),
  2195 => (x"7f",x"00",x"00",x"40"),
  2196 => (x"7f",x"19",x"09",x"7f"),
  2197 => (x"26",x"00",x"00",x"66"),
  2198 => (x"7b",x"59",x"4d",x"6f"),
  2199 => (x"01",x"00",x"00",x"32"),
  2200 => (x"01",x"7f",x"7f",x"01"),
  2201 => (x"3f",x"00",x"00",x"01"),
  2202 => (x"7f",x"40",x"40",x"7f"),
  2203 => (x"0f",x"00",x"00",x"3f"),
  2204 => (x"3f",x"70",x"70",x"3f"),
  2205 => (x"7f",x"7f",x"00",x"0f"),
  2206 => (x"7f",x"30",x"18",x"30"),
  2207 => (x"63",x"41",x"00",x"7f"),
  2208 => (x"36",x"1c",x"1c",x"36"),
  2209 => (x"03",x"01",x"41",x"63"),
  2210 => (x"06",x"7c",x"7c",x"06"),
  2211 => (x"71",x"61",x"01",x"03"),
  2212 => (x"43",x"47",x"4d",x"59"),
  2213 => (x"00",x"00",x"00",x"41"),
  2214 => (x"41",x"41",x"7f",x"7f"),
  2215 => (x"03",x"01",x"00",x"00"),
  2216 => (x"30",x"18",x"0c",x"06"),
  2217 => (x"00",x"00",x"40",x"60"),
  2218 => (x"7f",x"7f",x"41",x"41"),
  2219 => (x"0c",x"08",x"00",x"00"),
  2220 => (x"0c",x"06",x"03",x"06"),
  2221 => (x"80",x"80",x"00",x"08"),
  2222 => (x"80",x"80",x"80",x"80"),
  2223 => (x"00",x"00",x"00",x"80"),
  2224 => (x"04",x"07",x"03",x"00"),
  2225 => (x"20",x"00",x"00",x"00"),
  2226 => (x"7c",x"54",x"54",x"74"),
  2227 => (x"7f",x"00",x"00",x"78"),
  2228 => (x"7c",x"44",x"44",x"7f"),
  2229 => (x"38",x"00",x"00",x"38"),
  2230 => (x"44",x"44",x"44",x"7c"),
  2231 => (x"38",x"00",x"00",x"00"),
  2232 => (x"7f",x"44",x"44",x"7c"),
  2233 => (x"38",x"00",x"00",x"7f"),
  2234 => (x"5c",x"54",x"54",x"7c"),
  2235 => (x"04",x"00",x"00",x"18"),
  2236 => (x"05",x"05",x"7f",x"7e"),
  2237 => (x"18",x"00",x"00",x"00"),
  2238 => (x"fc",x"a4",x"a4",x"bc"),
  2239 => (x"7f",x"00",x"00",x"7c"),
  2240 => (x"7c",x"04",x"04",x"7f"),
  2241 => (x"00",x"00",x"00",x"78"),
  2242 => (x"40",x"7d",x"3d",x"00"),
  2243 => (x"80",x"00",x"00",x"00"),
  2244 => (x"7d",x"fd",x"80",x"80"),
  2245 => (x"7f",x"00",x"00",x"00"),
  2246 => (x"6c",x"38",x"10",x"7f"),
  2247 => (x"00",x"00",x"00",x"44"),
  2248 => (x"40",x"7f",x"3f",x"00"),
  2249 => (x"7c",x"7c",x"00",x"00"),
  2250 => (x"7c",x"0c",x"18",x"0c"),
  2251 => (x"7c",x"00",x"00",x"78"),
  2252 => (x"7c",x"04",x"04",x"7c"),
  2253 => (x"38",x"00",x"00",x"78"),
  2254 => (x"7c",x"44",x"44",x"7c"),
  2255 => (x"fc",x"00",x"00",x"38"),
  2256 => (x"3c",x"24",x"24",x"fc"),
  2257 => (x"18",x"00",x"00",x"18"),
  2258 => (x"fc",x"24",x"24",x"3c"),
  2259 => (x"7c",x"00",x"00",x"fc"),
  2260 => (x"0c",x"04",x"04",x"7c"),
  2261 => (x"48",x"00",x"00",x"08"),
  2262 => (x"74",x"54",x"54",x"5c"),
  2263 => (x"04",x"00",x"00",x"20"),
  2264 => (x"44",x"44",x"7f",x"3f"),
  2265 => (x"3c",x"00",x"00",x"00"),
  2266 => (x"7c",x"40",x"40",x"7c"),
  2267 => (x"1c",x"00",x"00",x"7c"),
  2268 => (x"3c",x"60",x"60",x"3c"),
  2269 => (x"7c",x"3c",x"00",x"1c"),
  2270 => (x"7c",x"60",x"30",x"60"),
  2271 => (x"6c",x"44",x"00",x"3c"),
  2272 => (x"6c",x"38",x"10",x"38"),
  2273 => (x"1c",x"00",x"00",x"44"),
  2274 => (x"3c",x"60",x"e0",x"bc"),
  2275 => (x"44",x"00",x"00",x"1c"),
  2276 => (x"4c",x"5c",x"74",x"64"),
  2277 => (x"08",x"00",x"00",x"44"),
  2278 => (x"41",x"77",x"3e",x"08"),
  2279 => (x"00",x"00",x"00",x"41"),
  2280 => (x"00",x"7f",x"7f",x"00"),
  2281 => (x"41",x"00",x"00",x"00"),
  2282 => (x"08",x"3e",x"77",x"41"),
  2283 => (x"01",x"02",x"00",x"08"),
  2284 => (x"02",x"02",x"03",x"01"),
  2285 => (x"7f",x"7f",x"00",x"01"),
  2286 => (x"7f",x"7f",x"7f",x"7f"),
  2287 => (x"08",x"08",x"00",x"7f"),
  2288 => (x"3e",x"3e",x"1c",x"1c"),
  2289 => (x"7f",x"7f",x"7f",x"7f"),
  2290 => (x"1c",x"1c",x"3e",x"3e"),
  2291 => (x"10",x"00",x"08",x"08"),
  2292 => (x"18",x"7c",x"7c",x"18"),
  2293 => (x"10",x"00",x"00",x"10"),
  2294 => (x"30",x"7c",x"7c",x"30"),
  2295 => (x"30",x"10",x"00",x"10"),
  2296 => (x"1e",x"78",x"60",x"60"),
  2297 => (x"66",x"42",x"00",x"06"),
  2298 => (x"66",x"3c",x"18",x"3c"),
  2299 => (x"38",x"78",x"00",x"42"),
  2300 => (x"6c",x"c6",x"c2",x"6a"),
  2301 => (x"00",x"60",x"00",x"38"),
  2302 => (x"00",x"00",x"60",x"00"),
  2303 => (x"5e",x"0e",x"00",x"60"),
  2304 => (x"0e",x"5d",x"5c",x"5b"),
  2305 => (x"c4",x"4c",x"71",x"1e"),
  2306 => (x"4d",x"bf",x"c2",x"cb"),
  2307 => (x"1e",x"c0",x"4b",x"c0"),
  2308 => (x"c7",x"02",x"ab",x"74"),
  2309 => (x"48",x"a6",x"c4",x"87"),
  2310 => (x"87",x"c5",x"78",x"c0"),
  2311 => (x"c1",x"48",x"a6",x"c4"),
  2312 => (x"1e",x"66",x"c4",x"78"),
  2313 => (x"df",x"ee",x"49",x"73"),
  2314 => (x"c0",x"86",x"c8",x"87"),
  2315 => (x"ef",x"ef",x"49",x"e0"),
  2316 => (x"4a",x"a5",x"c4",x"87"),
  2317 => (x"f0",x"f0",x"49",x"6a"),
  2318 => (x"87",x"c6",x"f1",x"87"),
  2319 => (x"83",x"c1",x"85",x"cb"),
  2320 => (x"04",x"ab",x"b7",x"c8"),
  2321 => (x"26",x"87",x"c7",x"ff"),
  2322 => (x"4c",x"26",x"4d",x"26"),
  2323 => (x"4f",x"26",x"4b",x"26"),
  2324 => (x"c4",x"4a",x"71",x"1e"),
  2325 => (x"c4",x"5a",x"c6",x"cb"),
  2326 => (x"c7",x"48",x"c6",x"cb"),
  2327 => (x"dd",x"fe",x"49",x"78"),
  2328 => (x"1e",x"4f",x"26",x"87"),
  2329 => (x"4a",x"71",x"1e",x"73"),
  2330 => (x"03",x"aa",x"b7",x"c0"),
  2331 => (x"df",x"c2",x"87",x"d3"),
  2332 => (x"c4",x"05",x"bf",x"f7"),
  2333 => (x"c2",x"4b",x"c1",x"87"),
  2334 => (x"c2",x"4b",x"c0",x"87"),
  2335 => (x"c4",x"5b",x"fb",x"df"),
  2336 => (x"fb",x"df",x"c2",x"87"),
  2337 => (x"f7",x"df",x"c2",x"5a"),
  2338 => (x"9a",x"c1",x"4a",x"bf"),
  2339 => (x"49",x"a2",x"c0",x"c1"),
  2340 => (x"fc",x"87",x"e8",x"ec"),
  2341 => (x"f7",x"df",x"c2",x"48"),
  2342 => (x"ef",x"fe",x"78",x"bf"),
  2343 => (x"4a",x"71",x"1e",x"87"),
  2344 => (x"72",x"1e",x"66",x"c4"),
  2345 => (x"87",x"f5",x"e9",x"49"),
  2346 => (x"1e",x"4f",x"26",x"26"),
  2347 => (x"bf",x"f7",x"df",x"c2"),
  2348 => (x"87",x"c8",x"e6",x"49"),
  2349 => (x"48",x"fa",x"ca",x"c4"),
  2350 => (x"c4",x"78",x"bf",x"e8"),
  2351 => (x"ec",x"48",x"f6",x"ca"),
  2352 => (x"ca",x"c4",x"78",x"bf"),
  2353 => (x"49",x"4a",x"bf",x"fa"),
  2354 => (x"ca",x"99",x"ff",x"cf"),
  2355 => (x"48",x"72",x"2a",x"b7"),
  2356 => (x"cb",x"c4",x"b0",x"71"),
  2357 => (x"4f",x"26",x"58",x"c2"),
  2358 => (x"5c",x"5b",x"5e",x"0e"),
  2359 => (x"4b",x"71",x"0e",x"5d"),
  2360 => (x"c4",x"87",x"c8",x"ff"),
  2361 => (x"c0",x"48",x"f5",x"ca"),
  2362 => (x"e5",x"49",x"73",x"50"),
  2363 => (x"49",x"70",x"87",x"f5"),
  2364 => (x"cb",x"9c",x"c2",x"4c"),
  2365 => (x"d7",x"c1",x"49",x"ee"),
  2366 => (x"49",x"70",x"87",x"cf"),
  2367 => (x"f5",x"ca",x"c4",x"4d"),
  2368 => (x"c1",x"05",x"bf",x"97"),
  2369 => (x"66",x"d0",x"87",x"e3"),
  2370 => (x"fe",x"ca",x"c4",x"49"),
  2371 => (x"d6",x"05",x"99",x"bf"),
  2372 => (x"49",x"66",x"d4",x"87"),
  2373 => (x"bf",x"f6",x"ca",x"c4"),
  2374 => (x"87",x"cb",x"05",x"99"),
  2375 => (x"c2",x"e5",x"49",x"73"),
  2376 => (x"02",x"98",x"70",x"87"),
  2377 => (x"c1",x"87",x"c2",x"c1"),
  2378 => (x"87",x"ff",x"fd",x"4c"),
  2379 => (x"d6",x"c1",x"49",x"75"),
  2380 => (x"98",x"70",x"87",x"e3"),
  2381 => (x"c4",x"87",x"c6",x"02"),
  2382 => (x"c1",x"48",x"f5",x"ca"),
  2383 => (x"f5",x"ca",x"c4",x"50"),
  2384 => (x"c0",x"05",x"bf",x"97"),
  2385 => (x"ca",x"c4",x"87",x"e3"),
  2386 => (x"d0",x"49",x"bf",x"fe"),
  2387 => (x"ff",x"05",x"99",x"66"),
  2388 => (x"ca",x"c4",x"87",x"d5"),
  2389 => (x"d4",x"49",x"bf",x"f6"),
  2390 => (x"ff",x"05",x"99",x"66"),
  2391 => (x"49",x"73",x"87",x"c9"),
  2392 => (x"70",x"87",x"c0",x"e4"),
  2393 => (x"fe",x"fe",x"05",x"98"),
  2394 => (x"fb",x"48",x"74",x"87"),
  2395 => (x"5e",x"0e",x"87",x"da"),
  2396 => (x"0e",x"5d",x"5c",x"5b"),
  2397 => (x"4d",x"c0",x"86",x"f4"),
  2398 => (x"7e",x"bf",x"ec",x"4c"),
  2399 => (x"c4",x"48",x"a6",x"c4"),
  2400 => (x"78",x"bf",x"c2",x"cb"),
  2401 => (x"1e",x"c0",x"1e",x"c1"),
  2402 => (x"cb",x"fd",x"49",x"c7"),
  2403 => (x"70",x"86",x"c8",x"87"),
  2404 => (x"87",x"cd",x"02",x"98"),
  2405 => (x"ca",x"fb",x"49",x"ff"),
  2406 => (x"49",x"da",x"c1",x"87"),
  2407 => (x"c1",x"87",x"c4",x"e3"),
  2408 => (x"f5",x"ca",x"c4",x"4d"),
  2409 => (x"c4",x"02",x"bf",x"97"),
  2410 => (x"ff",x"e0",x"c1",x"87"),
  2411 => (x"fa",x"ca",x"c4",x"87"),
  2412 => (x"df",x"c2",x"4b",x"bf"),
  2413 => (x"c1",x"05",x"bf",x"f7"),
  2414 => (x"a6",x"c4",x"87",x"da"),
  2415 => (x"c0",x"c0",x"c2",x"48"),
  2416 => (x"f8",x"c3",x"78",x"c0"),
  2417 => (x"97",x"6e",x"7e",x"fe"),
  2418 => (x"48",x"6e",x"49",x"bf"),
  2419 => (x"7e",x"70",x"80",x"c1"),
  2420 => (x"87",x"cf",x"e2",x"71"),
  2421 => (x"c3",x"02",x"98",x"70"),
  2422 => (x"b3",x"66",x"c4",x"87"),
  2423 => (x"c1",x"48",x"66",x"c4"),
  2424 => (x"a6",x"c8",x"28",x"b7"),
  2425 => (x"05",x"98",x"70",x"58"),
  2426 => (x"c3",x"87",x"db",x"ff"),
  2427 => (x"f2",x"e1",x"49",x"fd"),
  2428 => (x"49",x"fa",x"c3",x"87"),
  2429 => (x"73",x"87",x"ec",x"e1"),
  2430 => (x"99",x"ff",x"cf",x"49"),
  2431 => (x"49",x"c0",x"1e",x"71"),
  2432 => (x"73",x"87",x"da",x"fa"),
  2433 => (x"29",x"b7",x"ca",x"49"),
  2434 => (x"49",x"c1",x"1e",x"71"),
  2435 => (x"c8",x"87",x"ce",x"fa"),
  2436 => (x"87",x"c7",x"c6",x"86"),
  2437 => (x"bf",x"fe",x"ca",x"c4"),
  2438 => (x"df",x"02",x"9b",x"4b"),
  2439 => (x"f3",x"df",x"c2",x"87"),
  2440 => (x"d2",x"c1",x"49",x"bf"),
  2441 => (x"98",x"70",x"87",x"ef"),
  2442 => (x"c0",x"87",x"c4",x"05"),
  2443 => (x"c2",x"87",x"d3",x"4b"),
  2444 => (x"d2",x"c1",x"49",x"e0"),
  2445 => (x"df",x"c2",x"87",x"d3"),
  2446 => (x"87",x"c6",x"58",x"f7"),
  2447 => (x"48",x"f3",x"df",x"c2"),
  2448 => (x"49",x"73",x"78",x"c0"),
  2449 => (x"ce",x"05",x"99",x"c2"),
  2450 => (x"49",x"eb",x"c3",x"87"),
  2451 => (x"70",x"87",x"d4",x"e0"),
  2452 => (x"02",x"99",x"c2",x"49"),
  2453 => (x"fb",x"87",x"c2",x"c0"),
  2454 => (x"c1",x"49",x"73",x"4c"),
  2455 => (x"87",x"cf",x"05",x"99"),
  2456 => (x"ff",x"49",x"f4",x"c3"),
  2457 => (x"70",x"87",x"fc",x"df"),
  2458 => (x"02",x"99",x"c2",x"49"),
  2459 => (x"fa",x"87",x"c2",x"c0"),
  2460 => (x"c8",x"49",x"73",x"4c"),
  2461 => (x"87",x"ce",x"05",x"99"),
  2462 => (x"ff",x"49",x"f5",x"c3"),
  2463 => (x"70",x"87",x"e4",x"df"),
  2464 => (x"02",x"99",x"c2",x"49"),
  2465 => (x"cb",x"c4",x"87",x"d6"),
  2466 => (x"c0",x"02",x"bf",x"c6"),
  2467 => (x"c1",x"48",x"87",x"ca"),
  2468 => (x"ca",x"cb",x"c4",x"88"),
  2469 => (x"87",x"c2",x"c0",x"58"),
  2470 => (x"4d",x"c1",x"4c",x"ff"),
  2471 => (x"99",x"c4",x"49",x"73"),
  2472 => (x"87",x"ce",x"c0",x"05"),
  2473 => (x"ff",x"49",x"f2",x"c3"),
  2474 => (x"70",x"87",x"f8",x"de"),
  2475 => (x"02",x"99",x"c2",x"49"),
  2476 => (x"cb",x"c4",x"87",x"dc"),
  2477 => (x"48",x"7e",x"bf",x"c6"),
  2478 => (x"03",x"a8",x"b7",x"c7"),
  2479 => (x"6e",x"87",x"cb",x"c0"),
  2480 => (x"c4",x"80",x"c1",x"48"),
  2481 => (x"c0",x"58",x"ca",x"cb"),
  2482 => (x"4c",x"fe",x"87",x"c2"),
  2483 => (x"fd",x"c3",x"4d",x"c1"),
  2484 => (x"ce",x"de",x"ff",x"49"),
  2485 => (x"c2",x"49",x"70",x"87"),
  2486 => (x"d5",x"c0",x"02",x"99"),
  2487 => (x"c6",x"cb",x"c4",x"87"),
  2488 => (x"c9",x"c0",x"02",x"bf"),
  2489 => (x"c6",x"cb",x"c4",x"87"),
  2490 => (x"c0",x"78",x"c0",x"48"),
  2491 => (x"4c",x"fd",x"87",x"c2"),
  2492 => (x"fa",x"c3",x"4d",x"c1"),
  2493 => (x"ea",x"dd",x"ff",x"49"),
  2494 => (x"c2",x"49",x"70",x"87"),
  2495 => (x"d9",x"c0",x"02",x"99"),
  2496 => (x"c6",x"cb",x"c4",x"87"),
  2497 => (x"b7",x"c7",x"48",x"bf"),
  2498 => (x"c9",x"c0",x"03",x"a8"),
  2499 => (x"c6",x"cb",x"c4",x"87"),
  2500 => (x"c0",x"78",x"c7",x"48"),
  2501 => (x"4c",x"fc",x"87",x"c2"),
  2502 => (x"b7",x"c0",x"4d",x"c1"),
  2503 => (x"d1",x"c0",x"03",x"ac"),
  2504 => (x"4a",x"66",x"c4",x"87"),
  2505 => (x"6a",x"82",x"d8",x"c1"),
  2506 => (x"87",x"c6",x"c0",x"02"),
  2507 => (x"49",x"74",x"4b",x"6a"),
  2508 => (x"1e",x"c0",x"0f",x"73"),
  2509 => (x"c1",x"1e",x"f0",x"c3"),
  2510 => (x"db",x"f6",x"49",x"da"),
  2511 => (x"70",x"86",x"c8",x"87"),
  2512 => (x"e2",x"c0",x"02",x"98"),
  2513 => (x"48",x"a6",x"c8",x"87"),
  2514 => (x"bf",x"c6",x"cb",x"c4"),
  2515 => (x"49",x"66",x"c8",x"78"),
  2516 => (x"66",x"c4",x"91",x"cb"),
  2517 => (x"70",x"80",x"71",x"48"),
  2518 => (x"02",x"bf",x"6e",x"7e"),
  2519 => (x"6e",x"87",x"c8",x"c0"),
  2520 => (x"66",x"c8",x"4b",x"bf"),
  2521 => (x"75",x"0f",x"73",x"49"),
  2522 => (x"c8",x"c0",x"02",x"9d"),
  2523 => (x"c6",x"cb",x"c4",x"87"),
  2524 => (x"c9",x"f2",x"49",x"bf"),
  2525 => (x"fb",x"df",x"c2",x"87"),
  2526 => (x"de",x"c0",x"02",x"bf"),
  2527 => (x"cd",x"c1",x"49",x"87"),
  2528 => (x"98",x"70",x"87",x"d3"),
  2529 => (x"87",x"d3",x"c0",x"02"),
  2530 => (x"bf",x"c6",x"cb",x"c4"),
  2531 => (x"87",x"ee",x"f1",x"49"),
  2532 => (x"ce",x"f3",x"49",x"c0"),
  2533 => (x"fb",x"df",x"c2",x"87"),
  2534 => (x"f4",x"78",x"c0",x"48"),
  2535 => (x"87",x"e8",x"f2",x"8e"),
  2536 => (x"5c",x"5b",x"5e",x"0e"),
  2537 => (x"71",x"1e",x"0e",x"5d"),
  2538 => (x"c2",x"cb",x"c4",x"4c"),
  2539 => (x"cd",x"c1",x"49",x"bf"),
  2540 => (x"d1",x"c1",x"4d",x"a1"),
  2541 => (x"74",x"7e",x"69",x"81"),
  2542 => (x"87",x"cf",x"02",x"9c"),
  2543 => (x"74",x"4b",x"a5",x"c4"),
  2544 => (x"c2",x"cb",x"c4",x"7b"),
  2545 => (x"c7",x"f2",x"49",x"bf"),
  2546 => (x"74",x"7b",x"6e",x"87"),
  2547 => (x"87",x"c4",x"05",x"9c"),
  2548 => (x"87",x"c2",x"4b",x"c0"),
  2549 => (x"49",x"73",x"4b",x"c1"),
  2550 => (x"d4",x"87",x"c8",x"f2"),
  2551 => (x"87",x"c9",x"02",x"66"),
  2552 => (x"e4",x"cb",x"c1",x"49"),
  2553 => (x"c2",x"4a",x"70",x"87"),
  2554 => (x"c2",x"4a",x"c0",x"87"),
  2555 => (x"26",x"5a",x"ff",x"df"),
  2556 => (x"00",x"87",x"d5",x"f1"),
  2557 => (x"00",x"00",x"00",x"00"),
  2558 => (x"00",x"00",x"00",x"00"),
  2559 => (x"1e",x"00",x"00",x"00"),
  2560 => (x"4b",x"71",x"1e",x"73"),
  2561 => (x"4a",x"cb",x"c1",x"49"),
  2562 => (x"87",x"c7",x"e9",x"fd"),
  2563 => (x"72",x"1e",x"4a",x"70"),
  2564 => (x"4a",x"fc",x"c0",x"49"),
  2565 => (x"87",x"fb",x"e8",x"fd"),
  2566 => (x"4a",x"26",x"49",x"70"),
  2567 => (x"71",x"48",x"66",x"c8"),
  2568 => (x"c0",x"49",x"72",x"50"),
  2569 => (x"e8",x"fd",x"4a",x"fc"),
  2570 => (x"4a",x"71",x"87",x"e9"),
  2571 => (x"c1",x"49",x"66",x"c8"),
  2572 => (x"73",x"51",x"72",x"81"),
  2573 => (x"4a",x"cb",x"c1",x"49"),
  2574 => (x"87",x"d7",x"e8",x"fd"),
  2575 => (x"66",x"c8",x"4a",x"71"),
  2576 => (x"72",x"81",x"c2",x"49"),
  2577 => (x"26",x"87",x"c4",x"51"),
  2578 => (x"26",x"4c",x"26",x"4d"),
  2579 => (x"1e",x"4f",x"26",x"4b"),
  2580 => (x"4b",x"71",x"1e",x"73"),
  2581 => (x"c1",x"49",x"66",x"c8"),
  2582 => (x"66",x"cc",x"91",x"cb"),
  2583 => (x"73",x"49",x"a1",x"4a"),
  2584 => (x"d4",x"c6",x"c1",x"4a"),
  2585 => (x"49",x"a1",x"72",x"92"),
  2586 => (x"71",x"89",x"d6",x"c2"),
  2587 => (x"87",x"db",x"ff",x"48"),
  2588 => (x"5c",x"5b",x"5e",x"0e"),
  2589 => (x"71",x"1e",x"0e",x"5d"),
  2590 => (x"02",x"6b",x"97",x"4b"),
  2591 => (x"97",x"87",x"e4",x"c0"),
  2592 => (x"c0",x"48",x"7e",x"6b"),
  2593 => (x"04",x"a8",x"b7",x"f0"),
  2594 => (x"48",x"6e",x"87",x"d9"),
  2595 => (x"a8",x"b7",x"f9",x"c0"),
  2596 => (x"c1",x"87",x"d0",x"01"),
  2597 => (x"c0",x"49",x"6e",x"83"),
  2598 => (x"91",x"ca",x"89",x"f0"),
  2599 => (x"71",x"48",x"66",x"d4"),
  2600 => (x"c0",x"87",x"c5",x"50"),
  2601 => (x"87",x"eb",x"c4",x"48"),
  2602 => (x"c0",x"02",x"6b",x"97"),
  2603 => (x"6b",x"97",x"87",x"e9"),
  2604 => (x"f0",x"c0",x"48",x"7e"),
  2605 => (x"de",x"04",x"a8",x"b7"),
  2606 => (x"c0",x"48",x"6e",x"87"),
  2607 => (x"01",x"a8",x"b7",x"f9"),
  2608 => (x"83",x"c1",x"87",x"d5"),
  2609 => (x"f0",x"c0",x"49",x"6e"),
  2610 => (x"97",x"66",x"d4",x"89"),
  2611 => (x"49",x"a1",x"4a",x"bf"),
  2612 => (x"71",x"48",x"66",x"d4"),
  2613 => (x"c0",x"87",x"c5",x"50"),
  2614 => (x"87",x"f7",x"c3",x"48"),
  2615 => (x"cd",x"02",x"6b",x"97"),
  2616 => (x"49",x"6b",x"97",x"87"),
  2617 => (x"05",x"a9",x"fa",x"c0"),
  2618 => (x"83",x"c1",x"87",x"c4"),
  2619 => (x"48",x"c0",x"87",x"c5"),
  2620 => (x"97",x"87",x"e0",x"c3"),
  2621 => (x"e7",x"c0",x"02",x"6b"),
  2622 => (x"7e",x"6b",x"97",x"87"),
  2623 => (x"b7",x"f0",x"c0",x"48"),
  2624 => (x"87",x"dc",x"04",x"a8"),
  2625 => (x"f9",x"c0",x"48",x"6e"),
  2626 => (x"d3",x"01",x"a8",x"b7"),
  2627 => (x"6e",x"83",x"c1",x"87"),
  2628 => (x"89",x"f0",x"c0",x"49"),
  2629 => (x"66",x"d4",x"91",x"ca"),
  2630 => (x"71",x"84",x"c1",x"4c"),
  2631 => (x"87",x"c5",x"7c",x"97"),
  2632 => (x"ee",x"c2",x"48",x"c0"),
  2633 => (x"02",x"6b",x"97",x"87"),
  2634 => (x"97",x"87",x"e4",x"c0"),
  2635 => (x"c0",x"48",x"7e",x"6b"),
  2636 => (x"04",x"a8",x"b7",x"f0"),
  2637 => (x"48",x"6e",x"87",x"d9"),
  2638 => (x"a8",x"b7",x"f9",x"c0"),
  2639 => (x"c1",x"87",x"d0",x"01"),
  2640 => (x"c0",x"49",x"6e",x"83"),
  2641 => (x"6c",x"97",x"89",x"f0"),
  2642 => (x"97",x"49",x"a1",x"4a"),
  2643 => (x"c0",x"87",x"c5",x"7c"),
  2644 => (x"87",x"ff",x"c1",x"48"),
  2645 => (x"cd",x"02",x"6b",x"97"),
  2646 => (x"49",x"6b",x"97",x"87"),
  2647 => (x"05",x"a9",x"fa",x"c0"),
  2648 => (x"83",x"c1",x"87",x"c4"),
  2649 => (x"48",x"c0",x"87",x"c5"),
  2650 => (x"97",x"87",x"e8",x"c1"),
  2651 => (x"e4",x"c0",x"02",x"6b"),
  2652 => (x"4a",x"6b",x"97",x"87"),
  2653 => (x"aa",x"b7",x"f0",x"c0"),
  2654 => (x"c0",x"87",x"da",x"04"),
  2655 => (x"01",x"aa",x"b7",x"f9"),
  2656 => (x"83",x"c1",x"87",x"d3"),
  2657 => (x"f0",x"c0",x"49",x"72"),
  2658 => (x"d4",x"91",x"ca",x"89"),
  2659 => (x"85",x"c2",x"4d",x"66"),
  2660 => (x"c5",x"7d",x"97",x"71"),
  2661 => (x"c0",x"48",x"c0",x"87"),
  2662 => (x"6b",x"97",x"87",x"f9"),
  2663 => (x"87",x"e4",x"c0",x"02"),
  2664 => (x"48",x"7e",x"6b",x"97"),
  2665 => (x"a8",x"b7",x"f0",x"c0"),
  2666 => (x"6e",x"87",x"d9",x"04"),
  2667 => (x"b7",x"f9",x"c0",x"48"),
  2668 => (x"87",x"d0",x"01",x"a8"),
  2669 => (x"49",x"6e",x"83",x"c1"),
  2670 => (x"97",x"89",x"f0",x"c0"),
  2671 => (x"49",x"a1",x"4a",x"6d"),
  2672 => (x"87",x"c4",x"7d",x"97"),
  2673 => (x"87",x"cb",x"48",x"c0"),
  2674 => (x"c4",x"02",x"6b",x"97"),
  2675 => (x"c2",x"48",x"c0",x"87"),
  2676 => (x"26",x"48",x"c1",x"87"),
  2677 => (x"0e",x"87",x"f0",x"f9"),
  2678 => (x"5d",x"5c",x"5b",x"5e"),
  2679 => (x"71",x"86",x"f8",x"0e"),
  2680 => (x"4b",x"4c",x"c0",x"4d"),
  2681 => (x"49",x"c2",x"cc",x"c4"),
  2682 => (x"87",x"ff",x"cb",x"fe"),
  2683 => (x"b7",x"c0",x"4a",x"70"),
  2684 => (x"f2",x"c2",x"04",x"aa"),
  2685 => (x"02",x"aa",x"ca",x"87"),
  2686 => (x"c0",x"87",x"ec",x"c2"),
  2687 => (x"cf",x"02",x"aa",x"e0"),
  2688 => (x"02",x"aa",x"c9",x"87"),
  2689 => (x"aa",x"cd",x"87",x"ca"),
  2690 => (x"ca",x"87",x"c5",x"02"),
  2691 => (x"87",x"c6",x"05",x"aa"),
  2692 => (x"c2",x"02",x"9c",x"74"),
  2693 => (x"e2",x"c0",x"87",x"d1"),
  2694 => (x"87",x"cc",x"05",x"aa"),
  2695 => (x"b9",x"c1",x"49",x"74"),
  2696 => (x"ff",x"c3",x"4c",x"71"),
  2697 => (x"87",x"fc",x"fe",x"9c"),
  2698 => (x"c1",x"05",x"9c",x"74"),
  2699 => (x"e1",x"c1",x"87",x"e7"),
  2700 => (x"c8",x"04",x"aa",x"b7"),
  2701 => (x"b7",x"fa",x"c1",x"87"),
  2702 => (x"d8",x"c1",x"06",x"aa"),
  2703 => (x"b7",x"c1",x"c1",x"87"),
  2704 => (x"87",x"c8",x"04",x"aa"),
  2705 => (x"aa",x"b7",x"da",x"c1"),
  2706 => (x"87",x"c9",x"c1",x"06"),
  2707 => (x"aa",x"b7",x"f0",x"c0"),
  2708 => (x"c0",x"87",x"c8",x"04"),
  2709 => (x"06",x"aa",x"b7",x"f9"),
  2710 => (x"c1",x"87",x"fa",x"c0"),
  2711 => (x"c0",x"02",x"aa",x"db"),
  2712 => (x"dd",x"c1",x"87",x"f3"),
  2713 => (x"ec",x"c0",x"02",x"aa"),
  2714 => (x"aa",x"ed",x"c0",x"87"),
  2715 => (x"87",x"e5",x"c0",x"02"),
  2716 => (x"02",x"aa",x"df",x"c1"),
  2717 => (x"ec",x"c0",x"87",x"df"),
  2718 => (x"87",x"d9",x"02",x"aa"),
  2719 => (x"02",x"aa",x"fd",x"c0"),
  2720 => (x"fe",x"c1",x"87",x"d3"),
  2721 => (x"87",x"cd",x"02",x"aa"),
  2722 => (x"02",x"aa",x"fa",x"c0"),
  2723 => (x"ef",x"c0",x"87",x"c7"),
  2724 => (x"cf",x"fd",x"05",x"aa"),
  2725 => (x"b7",x"ff",x"c0",x"87"),
  2726 => (x"c7",x"fd",x"03",x"ab"),
  2727 => (x"49",x"a3",x"75",x"87"),
  2728 => (x"51",x"72",x"83",x"c1"),
  2729 => (x"75",x"87",x"fd",x"fc"),
  2730 => (x"51",x"c0",x"49",x"a3"),
  2731 => (x"c4",x"03",x"aa",x"b7"),
  2732 => (x"df",x"7e",x"c4",x"87"),
  2733 => (x"05",x"9b",x"73",x"87"),
  2734 => (x"a6",x"c4",x"87",x"c7"),
  2735 => (x"d0",x"78",x"c3",x"48"),
  2736 => (x"02",x"9c",x"74",x"87"),
  2737 => (x"7e",x"c1",x"87",x"c4"),
  2738 => (x"7e",x"c0",x"87",x"c2"),
  2739 => (x"6e",x"48",x"a6",x"c4"),
  2740 => (x"7e",x"66",x"c4",x"78"),
  2741 => (x"8e",x"f8",x"48",x"6e"),
  2742 => (x"0e",x"87",x"ec",x"f5"),
  2743 => (x"5d",x"5c",x"5b",x"5e"),
  2744 => (x"c4",x"4d",x"71",x"0e"),
  2745 => (x"c0",x"4b",x"ca",x"cb"),
  2746 => (x"49",x"f8",x"c0",x"4a"),
  2747 => (x"87",x"e6",x"d7",x"fd"),
  2748 => (x"cc",x"c4",x"1e",x"75"),
  2749 => (x"fc",x"fd",x"49",x"c2"),
  2750 => (x"86",x"c4",x"87",x"d4"),
  2751 => (x"c5",x"05",x"98",x"70"),
  2752 => (x"c0",x"4c",x"c1",x"87"),
  2753 => (x"49",x"c1",x"87",x"ea"),
  2754 => (x"70",x"87",x"ea",x"c0"),
  2755 => (x"c9",x"05",x"9c",x"4c"),
  2756 => (x"ce",x"cb",x"c4",x"87"),
  2757 => (x"87",x"dd",x"49",x"bf"),
  2758 => (x"9c",x"74",x"4c",x"70"),
  2759 => (x"c4",x"87",x"cb",x"05"),
  2760 => (x"c4",x"48",x"ca",x"cb"),
  2761 => (x"78",x"bf",x"de",x"cb"),
  2762 => (x"cb",x"c4",x"87",x"c6"),
  2763 => (x"78",x"c0",x"48",x"ce"),
  2764 => (x"d2",x"f4",x"48",x"74"),
  2765 => (x"5b",x"5e",x"0e",x"87"),
  2766 => (x"ff",x"0e",x"5d",x"5c"),
  2767 => (x"4c",x"71",x"86",x"d4"),
  2768 => (x"c4",x"7e",x"97",x"c0"),
  2769 => (x"50",x"c0",x"48",x"a6"),
  2770 => (x"c0",x"50",x"80",x"c0"),
  2771 => (x"80",x"c0",x"50",x"80"),
  2772 => (x"80",x"c0",x"4d",x"50"),
  2773 => (x"c0",x"80",x"c4",x"78"),
  2774 => (x"c0",x"80",x"c4",x"78"),
  2775 => (x"c0",x"80",x"c4",x"78"),
  2776 => (x"ca",x"cc",x"c4",x"78"),
  2777 => (x"87",x"c5",x"05",x"bf"),
  2778 => (x"c3",x"d0",x"48",x"c1"),
  2779 => (x"c2",x"cc",x"c4",x"87"),
  2780 => (x"d0",x"78",x"c0",x"48"),
  2781 => (x"f4",x"78",x"c0",x"80"),
  2782 => (x"ce",x"cc",x"c4",x"80"),
  2783 => (x"c0",x"c3",x"78",x"bf"),
  2784 => (x"78",x"c0",x"48",x"e2"),
  2785 => (x"48",x"de",x"cb",x"c4"),
  2786 => (x"ff",x"c2",x"78",x"c0"),
  2787 => (x"c6",x"f9",x"49",x"e2"),
  2788 => (x"58",x"a6",x"dc",x"87"),
  2789 => (x"cd",x"02",x"a8",x"c3"),
  2790 => (x"6e",x"97",x"87",x"d0"),
  2791 => (x"d8",x"02",x"9b",x"4b"),
  2792 => (x"02",x"8b",x"c1",x"87"),
  2793 => (x"8b",x"87",x"f5",x"c1"),
  2794 => (x"87",x"e4",x"c3",x"02"),
  2795 => (x"c4",x"c7",x"02",x"8b"),
  2796 => (x"c8",x"02",x"8b",x"87"),
  2797 => (x"f1",x"cc",x"87",x"c3"),
  2798 => (x"48",x"a6",x"c4",x"87"),
  2799 => (x"ff",x"c2",x"50",x"c0"),
  2800 => (x"fe",x"c2",x"4a",x"e2"),
  2801 => (x"d2",x"fd",x"49",x"d2"),
  2802 => (x"98",x"70",x"87",x"c5"),
  2803 => (x"c1",x"87",x"c6",x"05"),
  2804 => (x"d5",x"cc",x"7e",x"97"),
  2805 => (x"e2",x"ff",x"c2",x"87"),
  2806 => (x"d7",x"fe",x"c2",x"4a"),
  2807 => (x"ee",x"d1",x"fd",x"49"),
  2808 => (x"05",x"98",x"70",x"87"),
  2809 => (x"97",x"c2",x"87",x"c6"),
  2810 => (x"87",x"fe",x"cb",x"7e"),
  2811 => (x"4a",x"e2",x"ff",x"c2"),
  2812 => (x"49",x"dd",x"fe",x"c2"),
  2813 => (x"87",x"d7",x"d1",x"fd"),
  2814 => (x"c0",x"05",x"98",x"70"),
  2815 => (x"97",x"c3",x"87",x"c6"),
  2816 => (x"87",x"e6",x"cb",x"7e"),
  2817 => (x"4a",x"e2",x"ff",x"c2"),
  2818 => (x"49",x"e4",x"fe",x"c2"),
  2819 => (x"87",x"ff",x"d0",x"fd"),
  2820 => (x"cb",x"05",x"98",x"70"),
  2821 => (x"97",x"c4",x"87",x"d4"),
  2822 => (x"87",x"ce",x"cb",x"7e"),
  2823 => (x"48",x"66",x"97",x"c4"),
  2824 => (x"58",x"a6",x"e0",x"c0"),
  2825 => (x"c1",x"05",x"98",x"70"),
  2826 => (x"a6",x"c8",x"87",x"cd"),
  2827 => (x"c7",x"78",x"c0",x"48"),
  2828 => (x"c1",x"05",x"66",x"97"),
  2829 => (x"cb",x"c4",x"87",x"cd"),
  2830 => (x"c0",x"02",x"bf",x"f6"),
  2831 => (x"80",x"ff",x"87",x"c7"),
  2832 => (x"fe",x"c0",x"50",x"c1"),
  2833 => (x"e2",x"ff",x"c2",x"87"),
  2834 => (x"ee",x"cb",x"c4",x"1e"),
  2835 => (x"fd",x"f6",x"fd",x"49"),
  2836 => (x"70",x"86",x"c4",x"87"),
  2837 => (x"c8",x"c0",x"02",x"98"),
  2838 => (x"48",x"a6",x"c7",x"87"),
  2839 => (x"c5",x"c0",x"50",x"c1"),
  2840 => (x"48",x"a6",x"c5",x"87"),
  2841 => (x"f9",x"c3",x"50",x"c4"),
  2842 => (x"cc",x"c4",x"1e",x"fa"),
  2843 => (x"f9",x"fd",x"49",x"c2"),
  2844 => (x"86",x"c4",x"87",x"f8"),
  2845 => (x"dc",x"87",x"cc",x"c0"),
  2846 => (x"a8",x"c1",x"48",x"66"),
  2847 => (x"87",x"c3",x"c0",x"05"),
  2848 => (x"c4",x"7e",x"97",x"c0"),
  2849 => (x"c1",x"48",x"66",x"97"),
  2850 => (x"08",x"a6",x"c4",x"80"),
  2851 => (x"87",x"da",x"c9",x"50"),
  2852 => (x"c0",x"48",x"a6",x"d4"),
  2853 => (x"c4",x"78",x"66",x"e0"),
  2854 => (x"c0",x"48",x"66",x"97"),
  2855 => (x"70",x"58",x"a6",x"e0"),
  2856 => (x"fb",x"c0",x"05",x"98"),
  2857 => (x"c0",x"1e",x"ca",x"87"),
  2858 => (x"e2",x"ff",x"c2",x"1e"),
  2859 => (x"e0",x"d3",x"fd",x"49"),
  2860 => (x"70",x"86",x"c8",x"87"),
  2861 => (x"a6",x"e0",x"c0",x"49"),
  2862 => (x"02",x"66",x"dc",x"59"),
  2863 => (x"48",x"87",x"d3",x"c0"),
  2864 => (x"a8",x"b7",x"e3",x"c1"),
  2865 => (x"87",x"ca",x"c0",x"01"),
  2866 => (x"dc",x"49",x"a5",x"c1"),
  2867 => (x"c0",x"02",x"a9",x"66"),
  2868 => (x"a6",x"c5",x"87",x"c8"),
  2869 => (x"c2",x"50",x"c2",x"48"),
  2870 => (x"66",x"dc",x"87",x"ce"),
  2871 => (x"87",x"c8",x"c2",x"4d"),
  2872 => (x"c1",x"48",x"66",x"dc"),
  2873 => (x"ff",x"c1",x"05",x"a8"),
  2874 => (x"e2",x"ff",x"c2",x"87"),
  2875 => (x"f6",x"fd",x"c2",x"4a"),
  2876 => (x"da",x"cd",x"fd",x"49"),
  2877 => (x"05",x"98",x"70",x"87"),
  2878 => (x"c0",x"87",x"cf",x"c0"),
  2879 => (x"c0",x"48",x"a6",x"e0"),
  2880 => (x"c4",x"78",x"f0",x"e4"),
  2881 => (x"c1",x"78",x"c0",x"80"),
  2882 => (x"ff",x"c2",x"87",x"c7"),
  2883 => (x"fd",x"c2",x"4a",x"e2"),
  2884 => (x"cc",x"fd",x"49",x"fc"),
  2885 => (x"98",x"70",x"87",x"f9"),
  2886 => (x"87",x"cf",x"c0",x"05"),
  2887 => (x"48",x"a6",x"e0",x"c0"),
  2888 => (x"78",x"f0",x"e4",x"c0"),
  2889 => (x"78",x"c1",x"80",x"c4"),
  2890 => (x"c2",x"87",x"e6",x"c0"),
  2891 => (x"c2",x"4a",x"e2",x"ff"),
  2892 => (x"fd",x"49",x"c7",x"fe"),
  2893 => (x"70",x"87",x"d8",x"cc"),
  2894 => (x"cf",x"c0",x"05",x"98"),
  2895 => (x"a6",x"e0",x"c0",x"87"),
  2896 => (x"c0",x"e0",x"c0",x"48"),
  2897 => (x"c1",x"80",x"c4",x"78"),
  2898 => (x"87",x"c5",x"c0",x"78"),
  2899 => (x"c2",x"48",x"a6",x"c5"),
  2900 => (x"05",x"ac",x"75",x"50"),
  2901 => (x"c4",x"87",x"ce",x"c0"),
  2902 => (x"c0",x"48",x"e6",x"cb"),
  2903 => (x"fc",x"78",x"66",x"e0"),
  2904 => (x"66",x"e4",x"c0",x"80"),
  2905 => (x"7e",x"97",x"c0",x"78"),
  2906 => (x"48",x"66",x"97",x"c4"),
  2907 => (x"a6",x"c4",x"80",x"c1"),
  2908 => (x"f5",x"c5",x"50",x"08"),
  2909 => (x"a6",x"e8",x"c0",x"87"),
  2910 => (x"e2",x"ff",x"c2",x"1e"),
  2911 => (x"87",x"f0",x"eb",x"49"),
  2912 => (x"98",x"70",x"86",x"c4"),
  2913 => (x"87",x"c8",x"c0",x"05"),
  2914 => (x"c2",x"48",x"a6",x"c5"),
  2915 => (x"87",x"e3",x"c0",x"50"),
  2916 => (x"66",x"97",x"ea",x"c0"),
  2917 => (x"ed",x"c0",x"1e",x"49"),
  2918 => (x"1e",x"49",x"66",x"97"),
  2919 => (x"66",x"97",x"f0",x"c0"),
  2920 => (x"87",x"eb",x"ea",x"49"),
  2921 => (x"49",x"70",x"86",x"c8"),
  2922 => (x"71",x"81",x"d6",x"c2"),
  2923 => (x"80",x"66",x"c8",x"48"),
  2924 => (x"c0",x"58",x"a6",x"cc"),
  2925 => (x"f1",x"c4",x"7e",x"97"),
  2926 => (x"66",x"97",x"c4",x"87"),
  2927 => (x"a6",x"e0",x"c0",x"48"),
  2928 => (x"05",x"98",x"70",x"58"),
  2929 => (x"ca",x"87",x"d7",x"c0"),
  2930 => (x"c2",x"1e",x"c0",x"1e"),
  2931 => (x"fd",x"49",x"e2",x"ff"),
  2932 => (x"c8",x"87",x"fe",x"ce"),
  2933 => (x"ca",x"49",x"70",x"86"),
  2934 => (x"c4",x"59",x"97",x"a6"),
  2935 => (x"66",x"dc",x"87",x"c2"),
  2936 => (x"05",x"a8",x"c1",x"48"),
  2937 => (x"c0",x"87",x"f9",x"c3"),
  2938 => (x"c2",x"1e",x"a6",x"e8"),
  2939 => (x"e9",x"49",x"e2",x"ff"),
  2940 => (x"86",x"c4",x"87",x"fe"),
  2941 => (x"c0",x"05",x"98",x"70"),
  2942 => (x"a6",x"c5",x"87",x"c8"),
  2943 => (x"c3",x"50",x"c2",x"48"),
  2944 => (x"ea",x"c0",x"87",x"db"),
  2945 => (x"1e",x"49",x"66",x"97"),
  2946 => (x"66",x"97",x"ed",x"c0"),
  2947 => (x"f0",x"c0",x"1e",x"49"),
  2948 => (x"e8",x"49",x"66",x"97"),
  2949 => (x"86",x"c8",x"87",x"f9"),
  2950 => (x"97",x"c6",x"7e",x"70"),
  2951 => (x"e0",x"c0",x"48",x"66"),
  2952 => (x"98",x"70",x"58",x"a6"),
  2953 => (x"87",x"e1",x"c0",x"05"),
  2954 => (x"ad",x"49",x"a4",x"c1"),
  2955 => (x"87",x"ed",x"c2",x"05"),
  2956 => (x"bf",x"de",x"cb",x"c4"),
  2957 => (x"87",x"e5",x"c2",x"05"),
  2958 => (x"d6",x"c2",x"49",x"6e"),
  2959 => (x"c8",x"48",x"71",x"81"),
  2960 => (x"cb",x"c4",x"80",x"66"),
  2961 => (x"d4",x"c2",x"58",x"e2"),
  2962 => (x"48",x"66",x"dc",x"87"),
  2963 => (x"c2",x"05",x"a8",x"c1"),
  2964 => (x"ad",x"74",x"87",x"cb"),
  2965 => (x"87",x"ce",x"c0",x"05"),
  2966 => (x"d6",x"c2",x"49",x"6e"),
  2967 => (x"c8",x"48",x"71",x"81"),
  2968 => (x"cb",x"c4",x"80",x"66"),
  2969 => (x"b7",x"c1",x"58",x"de"),
  2970 => (x"ce",x"c1",x"06",x"ad"),
  2971 => (x"cc",x"48",x"6e",x"87"),
  2972 => (x"e0",x"c0",x"88",x"66"),
  2973 => (x"ad",x"74",x"58",x"a6"),
  2974 => (x"87",x"ce",x"c0",x"05"),
  2975 => (x"66",x"d4",x"49",x"70"),
  2976 => (x"d0",x"48",x"71",x"91"),
  2977 => (x"cb",x"c4",x"80",x"66"),
  2978 => (x"a4",x"c1",x"58",x"da"),
  2979 => (x"c0",x"05",x"ad",x"49"),
  2980 => (x"cb",x"c4",x"87",x"d8"),
  2981 => (x"c0",x"05",x"bf",x"de"),
  2982 => (x"49",x"6e",x"87",x"d0"),
  2983 => (x"c8",x"81",x"d6",x"c2"),
  2984 => (x"48",x"71",x"81",x"66"),
  2985 => (x"cb",x"c4",x"88",x"c1"),
  2986 => (x"66",x"dc",x"58",x"e2"),
  2987 => (x"91",x"66",x"d4",x"49"),
  2988 => (x"66",x"d0",x"48",x"71"),
  2989 => (x"58",x"a6",x"d4",x"80"),
  2990 => (x"6e",x"87",x"dd",x"c0"),
  2991 => (x"81",x"d6",x"c2",x"49"),
  2992 => (x"71",x"91",x"66",x"d4"),
  2993 => (x"80",x"66",x"d0",x"48"),
  2994 => (x"c1",x"58",x"a6",x"d4"),
  2995 => (x"c7",x"c0",x"05",x"ac"),
  2996 => (x"d6",x"cb",x"c4",x"87"),
  2997 => (x"78",x"66",x"d0",x"48"),
  2998 => (x"6e",x"48",x"a6",x"cc"),
  2999 => (x"7e",x"97",x"c0",x"78"),
  3000 => (x"48",x"66",x"97",x"c4"),
  3001 => (x"a6",x"c4",x"80",x"c1"),
  3002 => (x"66",x"d8",x"50",x"08"),
  3003 => (x"02",x"a8",x"c4",x"48"),
  3004 => (x"c5",x"87",x"c7",x"c0"),
  3005 => (x"f2",x"02",x"66",x"97"),
  3006 => (x"97",x"c7",x"87",x"d0"),
  3007 => (x"c8",x"c0",x"05",x"66"),
  3008 => (x"48",x"a6",x"c5",x"87"),
  3009 => (x"f1",x"c0",x"50",x"c4"),
  3010 => (x"05",x"ad",x"74",x"87"),
  3011 => (x"c4",x"87",x"eb",x"c0"),
  3012 => (x"4a",x"bf",x"d6",x"cb"),
  3013 => (x"bf",x"f6",x"cb",x"c4"),
  3014 => (x"70",x"88",x"72",x"48"),
  3015 => (x"e6",x"cb",x"c4",x"4a"),
  3016 => (x"1e",x"72",x"49",x"bf"),
  3017 => (x"fd",x"4a",x"09",x"72"),
  3018 => (x"70",x"87",x"f4",x"cb"),
  3019 => (x"c4",x"4a",x"26",x"49"),
  3020 => (x"48",x"bf",x"da",x"cb"),
  3021 => (x"cb",x"c4",x"80",x"71"),
  3022 => (x"b7",x"74",x"58",x"e2"),
  3023 => (x"c5",x"c0",x"03",x"ad"),
  3024 => (x"48",x"a6",x"c5",x"87"),
  3025 => (x"97",x"c5",x"50",x"c4"),
  3026 => (x"c9",x"c0",x"02",x"66"),
  3027 => (x"ce",x"cb",x"c4",x"87"),
  3028 => (x"c0",x"78",x"c0",x"48"),
  3029 => (x"cb",x"c4",x"87",x"c4"),
  3030 => (x"e8",x"c0",x"5d",x"d2"),
  3031 => (x"cb",x"c4",x"1e",x"a6"),
  3032 => (x"e2",x"49",x"bf",x"da"),
  3033 => (x"86",x"c4",x"87",x"d9"),
  3034 => (x"5c",x"ee",x"cb",x"c4"),
  3035 => (x"48",x"66",x"97",x"c5"),
  3036 => (x"e3",x"8e",x"d4",x"ff"),
  3037 => (x"55",x"41",x"87",x"d1"),
  3038 => (x"00",x"4f",x"49",x"44"),
  3039 => (x"45",x"44",x"4f",x"4d"),
  3040 => (x"33",x"32",x"2f",x"31"),
  3041 => (x"4d",x"00",x"32",x"35"),
  3042 => (x"31",x"45",x"44",x"4f"),
  3043 => (x"34",x"30",x"32",x"2f"),
  3044 => (x"49",x"46",x"00",x"38"),
  3045 => (x"54",x"00",x"45",x"4c"),
  3046 => (x"4b",x"43",x"41",x"52"),
  3047 => (x"45",x"52",x"50",x"00"),
  3048 => (x"00",x"50",x"41",x"47"),
  3049 => (x"45",x"44",x"4e",x"49"),
  3050 => (x"5e",x"0e",x"00",x"58"),
  3051 => (x"71",x"0e",x"5c",x"5b"),
  3052 => (x"c4",x"4c",x"c1",x"4b"),
  3053 => (x"b7",x"bf",x"da",x"cb"),
  3054 => (x"87",x"d0",x"04",x"ab"),
  3055 => (x"bf",x"de",x"cb",x"c4"),
  3056 => (x"c7",x"01",x"ab",x"b7"),
  3057 => (x"ea",x"cb",x"c4",x"87"),
  3058 => (x"87",x"d3",x"48",x"bf"),
  3059 => (x"e4",x"ed",x"49",x"74"),
  3060 => (x"c4",x"84",x"c1",x"87"),
  3061 => (x"b7",x"bf",x"ce",x"cb"),
  3062 => (x"d6",x"ff",x"06",x"ac"),
  3063 => (x"e1",x"48",x"ff",x"87"),
  3064 => (x"00",x"00",x"87",x"e7"),
  3065 => (x"00",x"00",x"00",x"00"),
  3066 => (x"00",x"00",x"00",x"00"),
  3067 => (x"00",x"00",x"00",x"00"),
  3068 => (x"00",x"00",x"00",x"00"),
  3069 => (x"00",x"00",x"00",x"00"),
  3070 => (x"00",x"00",x"00",x"00"),
  3071 => (x"00",x"00",x"00",x"00"),
  3072 => (x"00",x"00",x"00",x"00"),
  3073 => (x"00",x"00",x"00",x"00"),
  3074 => (x"00",x"00",x"00",x"00"),
  3075 => (x"00",x"00",x"00",x"00"),
  3076 => (x"00",x"00",x"00",x"00"),
  3077 => (x"00",x"00",x"00",x"00"),
  3078 => (x"00",x"00",x"00",x"00"),
  3079 => (x"00",x"00",x"00",x"00"),
  3080 => (x"00",x"00",x"00",x"00"),
  3081 => (x"73",x"1e",x"00",x"00"),
  3082 => (x"4a",x"4b",x"71",x"1e"),
  3083 => (x"ca",x"49",x"72",x"1e"),
  3084 => (x"de",x"c8",x"fd",x"4a"),
  3085 => (x"26",x"49",x"70",x"87"),
  3086 => (x"71",x"91",x"d0",x"4a"),
  3087 => (x"ca",x"49",x"72",x"1e"),
  3088 => (x"ce",x"c8",x"fd",x"4a"),
  3089 => (x"26",x"4a",x"71",x"87"),
  3090 => (x"49",x"a1",x"72",x"49"),
  3091 => (x"71",x"99",x"ff",x"c3"),
  3092 => (x"26",x"87",x"c4",x"48"),
  3093 => (x"26",x"4c",x"26",x"4d"),
  3094 => (x"1e",x"4f",x"26",x"4b"),
  3095 => (x"4b",x"71",x"1e",x"73"),
  3096 => (x"b7",x"c4",x"49",x"4a"),
  3097 => (x"cf",x"91",x"ca",x"29"),
  3098 => (x"49",x"a1",x"72",x"9a"),
  3099 => (x"71",x"99",x"ff",x"c3"),
  3100 => (x"1e",x"87",x"e4",x"48"),
  3101 => (x"4a",x"71",x"1e",x"73"),
  3102 => (x"70",x"87",x"e0",x"49"),
  3103 => (x"05",x"9b",x"4b",x"49"),
  3104 => (x"4b",x"c1",x"87",x"c2"),
  3105 => (x"bf",x"ce",x"cb",x"c4"),
  3106 => (x"c1",x"06",x"ab",x"b7"),
  3107 => (x"49",x"73",x"4b",x"87"),
  3108 => (x"73",x"87",x"e2",x"ea"),
  3109 => (x"87",x"ff",x"fe",x"48"),
  3110 => (x"ca",x"f1",x"c4",x"1e"),
  3111 => (x"f1",x"c4",x"59",x"97"),
  3112 => (x"66",x"c4",x"48",x"c7"),
  3113 => (x"50",x"66",x"c8",x"50"),
  3114 => (x"26",x"50",x"66",x"cc"),
  3115 => (x"1e",x"73",x"1e",x"4f"),
  3116 => (x"d0",x"ff",x"4b",x"71"),
  3117 => (x"78",x"c5",x"c8",x"48"),
  3118 => (x"c1",x"48",x"d4",x"ff"),
  3119 => (x"49",x"73",x"78",x"e1"),
  3120 => (x"2a",x"b7",x"c8",x"4a"),
  3121 => (x"ff",x"c3",x"78",x"72"),
  3122 => (x"ff",x"78",x"71",x"99"),
  3123 => (x"78",x"c4",x"48",x"d0"),
  3124 => (x"1e",x"87",x"c4",x"fe"),
  3125 => (x"9f",x"c4",x"f2",x"c4"),
  3126 => (x"d4",x"f1",x"c4",x"59"),
  3127 => (x"26",x"78",x"c1",x"48"),
  3128 => (x"5b",x"5e",x"0e",x"4f"),
  3129 => (x"4c",x"71",x"0e",x"5c"),
  3130 => (x"c8",x"48",x"d0",x"ff"),
  3131 => (x"d4",x"ff",x"78",x"c5"),
  3132 => (x"78",x"e4",x"c1",x"48"),
  3133 => (x"4a",x"49",x"66",x"cc"),
  3134 => (x"72",x"9a",x"ff",x"c3"),
  3135 => (x"4a",x"66",x"cc",x"78"),
  3136 => (x"ff",x"c3",x"2a",x"c8"),
  3137 => (x"4b",x"66",x"d0",x"9a"),
  3138 => (x"b2",x"73",x"33",x"c7"),
  3139 => (x"1e",x"71",x"78",x"72"),
  3140 => (x"c5",x"fd",x"49",x"74"),
  3141 => (x"d0",x"ff",x"87",x"ee"),
  3142 => (x"26",x"78",x"c4",x"48"),
  3143 => (x"1e",x"87",x"f6",x"fc"),
  3144 => (x"e0",x"c0",x"1e",x"73"),
  3145 => (x"cb",x"c4",x"4b",x"c0"),
  3146 => (x"c1",x"02",x"bf",x"e2"),
  3147 => (x"f1",x"c4",x"87",x"e7"),
  3148 => (x"c0",x"48",x"bf",x"df"),
  3149 => (x"c1",x"04",x"a8",x"b7"),
  3150 => (x"cb",x"c4",x"87",x"db"),
  3151 => (x"02",x"ab",x"bf",x"e6"),
  3152 => (x"cb",x"c4",x"87",x"d3"),
  3153 => (x"d0",x"49",x"bf",x"fe"),
  3154 => (x"c4",x"1e",x"71",x"81"),
  3155 => (x"fd",x"49",x"ee",x"cb"),
  3156 => (x"c4",x"87",x"dd",x"e8"),
  3157 => (x"c4",x"1e",x"73",x"86"),
  3158 => (x"c4",x"1e",x"d6",x"cc"),
  3159 => (x"fd",x"49",x"ee",x"cb"),
  3160 => (x"c8",x"87",x"f4",x"e9"),
  3161 => (x"e6",x"cb",x"c4",x"86"),
  3162 => (x"d6",x"02",x"ab",x"bf"),
  3163 => (x"e0",x"c0",x"49",x"87"),
  3164 => (x"cb",x"c4",x"89",x"d0"),
  3165 => (x"71",x"81",x"bf",x"fe"),
  3166 => (x"ee",x"cb",x"c4",x"1e"),
  3167 => (x"ef",x"e7",x"fd",x"49"),
  3168 => (x"c8",x"86",x"c4",x"87"),
  3169 => (x"73",x"1e",x"49",x"66"),
  3170 => (x"d6",x"cc",x"c4",x"1e"),
  3171 => (x"87",x"d1",x"fd",x"49"),
  3172 => (x"e1",x"c0",x"86",x"c8"),
  3173 => (x"f0",x"e4",x"c0",x"87"),
  3174 => (x"d6",x"cc",x"c4",x"1e"),
  3175 => (x"ee",x"cb",x"c4",x"1e"),
  3176 => (x"f2",x"e8",x"fd",x"49"),
  3177 => (x"49",x"66",x"d0",x"87"),
  3178 => (x"f0",x"e4",x"c0",x"1e"),
  3179 => (x"d6",x"cc",x"c4",x"1e"),
  3180 => (x"87",x"ed",x"fc",x"49"),
  3181 => (x"de",x"fa",x"86",x"d0"),
  3182 => (x"cb",x"c4",x"1e",x"87"),
  3183 => (x"db",x"05",x"bf",x"f6"),
  3184 => (x"ce",x"f1",x"c4",x"87"),
  3185 => (x"c0",x"50",x"c1",x"48"),
  3186 => (x"1e",x"cb",x"1e",x"1e"),
  3187 => (x"c7",x"fb",x"49",x"c2"),
  3188 => (x"c1",x"86",x"cc",x"87"),
  3189 => (x"87",x"d5",x"fb",x"49"),
  3190 => (x"87",x"c2",x"48",x"c0"),
  3191 => (x"4f",x"26",x"48",x"c1"),
  3192 => (x"c4",x"1e",x"73",x"1e"),
  3193 => (x"48",x"bf",x"ca",x"f1"),
  3194 => (x"c0",x"06",x"a8",x"c0"),
  3195 => (x"eb",x"c3",x"87",x"e9"),
  3196 => (x"c0",x"49",x"bf",x"c5"),
  3197 => (x"70",x"87",x"de",x"e3"),
  3198 => (x"e3",x"c7",x"02",x"98"),
  3199 => (x"c0",x"49",x"cd",x"87"),
  3200 => (x"70",x"87",x"c6",x"e3"),
  3201 => (x"c9",x"eb",x"c3",x"49"),
  3202 => (x"ca",x"f1",x"c4",x"59"),
  3203 => (x"88",x"c1",x"48",x"bf"),
  3204 => (x"58",x"ce",x"f1",x"c4"),
  3205 => (x"c4",x"87",x"c9",x"c7"),
  3206 => (x"bf",x"97",x"ce",x"f1"),
  3207 => (x"05",x"aa",x"c2",x"4a"),
  3208 => (x"c4",x"87",x"ca",x"c3"),
  3209 => (x"48",x"bf",x"db",x"f1"),
  3210 => (x"bf",x"ce",x"cb",x"c4"),
  3211 => (x"c9",x"06",x"a8",x"b7"),
  3212 => (x"ce",x"f1",x"c4",x"87"),
  3213 => (x"c6",x"50",x"c0",x"48"),
  3214 => (x"f1",x"c4",x"87",x"e6"),
  3215 => (x"02",x"bf",x"97",x"d9"),
  3216 => (x"c4",x"87",x"dd",x"c6"),
  3217 => (x"05",x"bf",x"f6",x"cb"),
  3218 => (x"f1",x"c4",x"87",x"da"),
  3219 => (x"50",x"c1",x"48",x"ce"),
  3220 => (x"cb",x"1e",x"1e",x"c0"),
  3221 => (x"f8",x"49",x"c2",x"1e"),
  3222 => (x"86",x"cc",x"87",x"fe"),
  3223 => (x"f2",x"f9",x"49",x"c1"),
  3224 => (x"87",x"fc",x"c5",x"87"),
  3225 => (x"48",x"d9",x"f1",x"c4"),
  3226 => (x"cb",x"c4",x"50",x"c0"),
  3227 => (x"cd",x"02",x"bf",x"e2"),
  3228 => (x"c0",x"1e",x"c1",x"87"),
  3229 => (x"fa",x"49",x"c0",x"e0"),
  3230 => (x"86",x"c4",x"87",x"e5"),
  3231 => (x"f1",x"c4",x"87",x"d5"),
  3232 => (x"c4",x"48",x"bf",x"df"),
  3233 => (x"b7",x"bf",x"da",x"cb"),
  3234 => (x"c6",x"c0",x"04",x"a8"),
  3235 => (x"cf",x"f1",x"c4",x"87"),
  3236 => (x"c4",x"50",x"c0",x"48"),
  3237 => (x"48",x"bf",x"e3",x"f1"),
  3238 => (x"f1",x"c4",x"88",x"c1"),
  3239 => (x"98",x"70",x"58",x"e7"),
  3240 => (x"87",x"cb",x"c0",x"05"),
  3241 => (x"ea",x"f8",x"49",x"c0"),
  3242 => (x"ce",x"f1",x"c4",x"87"),
  3243 => (x"c4",x"50",x"c0",x"48"),
  3244 => (x"48",x"bf",x"df",x"f1"),
  3245 => (x"f1",x"c4",x"80",x"c1"),
  3246 => (x"cb",x"c4",x"58",x"e3"),
  3247 => (x"a8",x"b7",x"bf",x"de"),
  3248 => (x"87",x"dc",x"c4",x"04"),
  3249 => (x"bf",x"db",x"f1",x"c4"),
  3250 => (x"c4",x"80",x"c1",x"48"),
  3251 => (x"70",x"58",x"df",x"f1"),
  3252 => (x"87",x"e1",x"e1",x"49"),
  3253 => (x"48",x"cf",x"f1",x"c4"),
  3254 => (x"cb",x"c4",x"50",x"c1"),
  3255 => (x"1e",x"49",x"bf",x"d6"),
  3256 => (x"49",x"ee",x"cb",x"c4"),
  3257 => (x"87",x"c8",x"e2",x"fd"),
  3258 => (x"f3",x"c3",x"86",x"c4"),
  3259 => (x"05",x"aa",x"c3",x"87"),
  3260 => (x"c4",x"87",x"ed",x"c3"),
  3261 => (x"05",x"bf",x"f6",x"cb"),
  3262 => (x"c4",x"87",x"da",x"c0"),
  3263 => (x"c1",x"48",x"ce",x"f1"),
  3264 => (x"1e",x"1e",x"c0",x"50"),
  3265 => (x"49",x"c2",x"1e",x"cb"),
  3266 => (x"cc",x"87",x"cd",x"f6"),
  3267 => (x"f7",x"49",x"c1",x"86"),
  3268 => (x"cb",x"c3",x"87",x"c1"),
  3269 => (x"df",x"f1",x"c4",x"87"),
  3270 => (x"cd",x"f2",x"49",x"bf"),
  3271 => (x"df",x"f1",x"c4",x"87"),
  3272 => (x"da",x"f1",x"c4",x"58"),
  3273 => (x"c1",x"05",x"bf",x"97"),
  3274 => (x"4b",x"c0",x"87",x"d5"),
  3275 => (x"bf",x"fb",x"f1",x"c4"),
  3276 => (x"a8",x"b7",x"c0",x"48"),
  3277 => (x"87",x"c7",x"c1",x"04"),
  3278 => (x"bf",x"e2",x"cb",x"c4"),
  3279 => (x"87",x"e8",x"c0",x"05"),
  3280 => (x"bf",x"df",x"f1",x"c4"),
  3281 => (x"da",x"cb",x"c4",x"49"),
  3282 => (x"e4",x"c0",x"89",x"bf"),
  3283 => (x"cb",x"c4",x"91",x"f0"),
  3284 => (x"71",x"81",x"bf",x"d6"),
  3285 => (x"ee",x"cb",x"c4",x"1e"),
  3286 => (x"d3",x"e0",x"fd",x"49"),
  3287 => (x"c0",x"1e",x"c0",x"87"),
  3288 => (x"f6",x"49",x"f0",x"e4"),
  3289 => (x"86",x"c8",x"87",x"f9"),
  3290 => (x"bf",x"df",x"f1",x"c4"),
  3291 => (x"c4",x"80",x"c1",x"48"),
  3292 => (x"c1",x"58",x"e3",x"f1"),
  3293 => (x"fb",x"f1",x"c4",x"83"),
  3294 => (x"06",x"ab",x"b7",x"bf"),
  3295 => (x"c4",x"87",x"f9",x"fe"),
  3296 => (x"c0",x"48",x"fb",x"f1"),
  3297 => (x"df",x"f1",x"c4",x"78"),
  3298 => (x"f1",x"c4",x"48",x"bf"),
  3299 => (x"a8",x"b7",x"bf",x"f7"),
  3300 => (x"87",x"d7",x"c0",x"03"),
  3301 => (x"bf",x"e2",x"cb",x"c4"),
  3302 => (x"87",x"cf",x"c0",x"05"),
  3303 => (x"bf",x"db",x"f1",x"c4"),
  3304 => (x"ce",x"cb",x"c4",x"48"),
  3305 => (x"06",x"a8",x"b7",x"bf"),
  3306 => (x"c4",x"87",x"f5",x"c0"),
  3307 => (x"bf",x"97",x"ff",x"f1"),
  3308 => (x"05",x"a9",x"c1",x"49"),
  3309 => (x"c4",x"87",x"d2",x"c0"),
  3310 => (x"c4",x"48",x"df",x"f1"),
  3311 => (x"78",x"bf",x"f3",x"f1"),
  3312 => (x"48",x"ca",x"f1",x"c4"),
  3313 => (x"c6",x"c0",x"78",x"c2"),
  3314 => (x"ce",x"f1",x"c4",x"87"),
  3315 => (x"c4",x"50",x"c0",x"48"),
  3316 => (x"bf",x"97",x"ff",x"f1"),
  3317 => (x"05",x"a9",x"c2",x"49"),
  3318 => (x"c0",x"87",x"c5",x"c0"),
  3319 => (x"87",x"f3",x"f3",x"49"),
  3320 => (x"0e",x"87",x"f4",x"f1"),
  3321 => (x"5d",x"5c",x"5b",x"5e"),
  3322 => (x"86",x"c4",x"ff",x"0e"),
  3323 => (x"4a",x"c0",x"4b",x"76"),
  3324 => (x"fc",x"49",x"e0",x"c0"),
  3325 => (x"ff",x"87",x"df",x"f3"),
  3326 => (x"c5",x"c8",x"48",x"d0"),
  3327 => (x"48",x"d4",x"ff",x"78"),
  3328 => (x"c0",x"78",x"e2",x"c1"),
  3329 => (x"c0",x"48",x"a6",x"e0"),
  3330 => (x"48",x"d4",x"ff",x"78"),
  3331 => (x"e4",x"c0",x"78",x"c0"),
  3332 => (x"e0",x"c0",x"49",x"a6"),
  3333 => (x"51",x"68",x"81",x"66"),
  3334 => (x"48",x"66",x"e0",x"c0"),
  3335 => (x"e4",x"c0",x"80",x"c1"),
  3336 => (x"b7",x"cc",x"58",x"a6"),
  3337 => (x"e0",x"ff",x"04",x"a8"),
  3338 => (x"48",x"d0",x"ff",x"87"),
  3339 => (x"e4",x"c0",x"78",x"c4"),
  3340 => (x"9c",x"4c",x"66",x"97"),
  3341 => (x"87",x"f3",x"c0",x"02"),
  3342 => (x"c0",x"02",x"8c",x"c3"),
  3343 => (x"8c",x"c5",x"87",x"fe"),
  3344 => (x"87",x"e5",x"c6",x"02"),
  3345 => (x"c8",x"02",x"8c",x"cd"),
  3346 => (x"c3",x"c3",x"87",x"e9"),
  3347 => (x"fb",x"c8",x"02",x"8c"),
  3348 => (x"02",x"8c",x"c1",x"87"),
  3349 => (x"8c",x"87",x"d2",x"cc"),
  3350 => (x"87",x"c9",x"d0",x"02"),
  3351 => (x"d0",x"02",x"8c",x"c3"),
  3352 => (x"8c",x"c1",x"87",x"da"),
  3353 => (x"87",x"f8",x"c1",x"02"),
  3354 => (x"f5",x"87",x"cc",x"d4"),
  3355 => (x"98",x"70",x"87",x"cb"),
  3356 => (x"87",x"dd",x"d4",x"02"),
  3357 => (x"f4",x"f0",x"49",x"c0"),
  3358 => (x"87",x"d5",x"d4",x"87"),
  3359 => (x"c1",x"7e",x"97",x"d2"),
  3360 => (x"c0",x"c2",x"48",x"a6"),
  3361 => (x"50",x"f0",x"c1",x"50"),
  3362 => (x"f1",x"c4",x"80",x"c1"),
  3363 => (x"50",x"bf",x"97",x"c6"),
  3364 => (x"50",x"ca",x"80",x"c4"),
  3365 => (x"f1",x"c4",x"80",x"c4"),
  3366 => (x"50",x"bf",x"97",x"c7"),
  3367 => (x"97",x"c8",x"f1",x"c4"),
  3368 => (x"f1",x"c4",x"50",x"bf"),
  3369 => (x"50",x"bf",x"97",x"c9"),
  3370 => (x"48",x"c9",x"f1",x"c4"),
  3371 => (x"f1",x"c4",x"50",x"c0"),
  3372 => (x"f1",x"c4",x"48",x"c8"),
  3373 => (x"50",x"bf",x"97",x"c9"),
  3374 => (x"48",x"c7",x"f1",x"c4"),
  3375 => (x"97",x"c8",x"f1",x"c4"),
  3376 => (x"f1",x"c4",x"50",x"bf"),
  3377 => (x"f1",x"c4",x"48",x"c6"),
  3378 => (x"50",x"bf",x"97",x"c7"),
  3379 => (x"1e",x"d2",x"1e",x"c1"),
  3380 => (x"f0",x"49",x"a6",x"ca"),
  3381 => (x"86",x"c8",x"87",x"cb"),
  3382 => (x"d0",x"ef",x"49",x"c0"),
  3383 => (x"87",x"f1",x"d2",x"87"),
  3384 => (x"70",x"87",x"d6",x"f3"),
  3385 => (x"e8",x"d2",x"02",x"98"),
  3386 => (x"97",x"e5",x"c0",x"87"),
  3387 => (x"e4",x"c0",x"48",x"66"),
  3388 => (x"98",x"70",x"58",x"a6"),
  3389 => (x"48",x"87",x"da",x"02"),
  3390 => (x"e4",x"c0",x"88",x"c1"),
  3391 => (x"98",x"70",x"58",x"a6"),
  3392 => (x"87",x"ed",x"c0",x"02"),
  3393 => (x"c0",x"88",x"c1",x"48"),
  3394 => (x"70",x"58",x"a6",x"e4"),
  3395 => (x"eb",x"c1",x"02",x"98"),
  3396 => (x"7e",x"97",x"c2",x"87"),
  3397 => (x"c2",x"48",x"a6",x"c1"),
  3398 => (x"50",x"c1",x"50",x"c0"),
  3399 => (x"bf",x"ce",x"cb",x"c4"),
  3400 => (x"87",x"c2",x"ec",x"49"),
  3401 => (x"50",x"08",x"a6",x"c3"),
  3402 => (x"48",x"a6",x"e0",x"c0"),
  3403 => (x"e2",x"c2",x"78",x"c2"),
  3404 => (x"ca",x"cb",x"c4",x"87"),
  3405 => (x"d6",x"c2",x"49",x"bf"),
  3406 => (x"a6",x"f0",x"c0",x"81"),
  3407 => (x"ca",x"ff",x"71",x"1e"),
  3408 => (x"86",x"c4",x"87",x"fd"),
  3409 => (x"a6",x"c1",x"7e",x"97"),
  3410 => (x"50",x"c0",x"c2",x"48"),
  3411 => (x"66",x"97",x"f0",x"c0"),
  3412 => (x"87",x"d2",x"eb",x"49"),
  3413 => (x"50",x"08",x"a6",x"c2"),
  3414 => (x"66",x"97",x"f1",x"c0"),
  3415 => (x"87",x"c6",x"eb",x"49"),
  3416 => (x"50",x"08",x"a6",x"c3"),
  3417 => (x"66",x"97",x"f2",x"c0"),
  3418 => (x"87",x"fa",x"ea",x"49"),
  3419 => (x"50",x"08",x"a6",x"c4"),
  3420 => (x"c0",x"48",x"a6",x"c5"),
  3421 => (x"c4",x"80",x"da",x"50"),
  3422 => (x"87",x"d7",x"c1",x"78"),
  3423 => (x"66",x"97",x"e6",x"c0"),
  3424 => (x"87",x"ef",x"eb",x"49"),
  3425 => (x"bf",x"da",x"cb",x"c4"),
  3426 => (x"81",x"d6",x"c2",x"49"),
  3427 => (x"1e",x"a6",x"f0",x"c0"),
  3428 => (x"ea",x"c9",x"ff",x"71"),
  3429 => (x"97",x"86",x"c4",x"87"),
  3430 => (x"48",x"a6",x"c1",x"7e"),
  3431 => (x"c0",x"50",x"c0",x"c2"),
  3432 => (x"49",x"66",x"97",x"f0"),
  3433 => (x"c2",x"87",x"ff",x"e9"),
  3434 => (x"c0",x"50",x"08",x"a6"),
  3435 => (x"49",x"66",x"97",x"f1"),
  3436 => (x"c3",x"87",x"f3",x"e9"),
  3437 => (x"c0",x"50",x"08",x"a6"),
  3438 => (x"49",x"66",x"97",x"f2"),
  3439 => (x"c4",x"87",x"e7",x"e9"),
  3440 => (x"c4",x"50",x"08",x"a6"),
  3441 => (x"49",x"bf",x"e2",x"cb"),
  3442 => (x"a6",x"c9",x"31",x"c2"),
  3443 => (x"db",x"48",x"59",x"97"),
  3444 => (x"c1",x"78",x"c4",x"80"),
  3445 => (x"66",x"e4",x"c0",x"1e"),
  3446 => (x"49",x"a6",x"ca",x"1e"),
  3447 => (x"c8",x"87",x"c2",x"ec"),
  3448 => (x"eb",x"49",x"c0",x"86"),
  3449 => (x"e8",x"ce",x"87",x"c7"),
  3450 => (x"87",x"cd",x"ef",x"87"),
  3451 => (x"ce",x"02",x"98",x"70"),
  3452 => (x"e5",x"c0",x"87",x"df"),
  3453 => (x"d0",x"49",x"66",x"97"),
  3454 => (x"97",x"e6",x"c0",x"31"),
  3455 => (x"32",x"c8",x"4a",x"66"),
  3456 => (x"e7",x"c0",x"b1",x"72"),
  3457 => (x"b1",x"4a",x"66",x"97"),
  3458 => (x"ff",x"c7",x"4d",x"71"),
  3459 => (x"c0",x"9d",x"ff",x"ff"),
  3460 => (x"02",x"66",x"97",x"e8"),
  3461 => (x"48",x"87",x"c8",x"c0"),
  3462 => (x"58",x"a6",x"e4",x"c0"),
  3463 => (x"c0",x"87",x"c7",x"c0"),
  3464 => (x"c4",x"48",x"a6",x"e0"),
  3465 => (x"49",x"75",x"78",x"c0"),
  3466 => (x"c4",x"87",x"ff",x"e5"),
  3467 => (x"c4",x"58",x"df",x"f1"),
  3468 => (x"c0",x"48",x"ca",x"f1"),
  3469 => (x"e3",x"f1",x"c4",x"78"),
  3470 => (x"e3",x"f1",x"c4",x"5d"),
  3471 => (x"66",x"e0",x"c0",x"48"),
  3472 => (x"c4",x"49",x"75",x"78"),
  3473 => (x"89",x"bf",x"da",x"cb"),
  3474 => (x"bf",x"e6",x"cb",x"c4"),
  3475 => (x"d6",x"cb",x"c4",x"91"),
  3476 => (x"1e",x"71",x"81",x"bf"),
  3477 => (x"49",x"ee",x"cb",x"c4"),
  3478 => (x"87",x"d4",x"d4",x"fd"),
  3479 => (x"f1",x"c4",x"86",x"c4"),
  3480 => (x"78",x"c0",x"48",x"ef"),
  3481 => (x"48",x"d9",x"f1",x"c4"),
  3482 => (x"f1",x"c4",x"50",x"c1"),
  3483 => (x"50",x"c2",x"48",x"ce"),
  3484 => (x"c0",x"87",x"de",x"cc"),
  3485 => (x"02",x"66",x"97",x"e8"),
  3486 => (x"c4",x"87",x"c9",x"c0"),
  3487 => (x"c1",x"48",x"d8",x"f1"),
  3488 => (x"87",x"cd",x"cc",x"50"),
  3489 => (x"e4",x"e8",x"49",x"c0"),
  3490 => (x"87",x"c5",x"cc",x"87"),
  3491 => (x"70",x"87",x"ea",x"ec"),
  3492 => (x"fc",x"cb",x"02",x"98"),
  3493 => (x"97",x"ed",x"c0",x"87"),
  3494 => (x"c3",x"48",x"49",x"66"),
  3495 => (x"e4",x"c0",x"98",x"c0"),
  3496 => (x"98",x"70",x"58",x"a6"),
  3497 => (x"87",x"dc",x"c0",x"02"),
  3498 => (x"88",x"c0",x"c1",x"48"),
  3499 => (x"58",x"a6",x"e4",x"c0"),
  3500 => (x"c0",x"02",x"98",x"70"),
  3501 => (x"c1",x"48",x"87",x"e9"),
  3502 => (x"e4",x"c0",x"88",x"c0"),
  3503 => (x"98",x"70",x"58",x"a6"),
  3504 => (x"87",x"c7",x"c1",x"02"),
  3505 => (x"66",x"97",x"e7",x"c0"),
  3506 => (x"c0",x"31",x"d0",x"49"),
  3507 => (x"4a",x"66",x"97",x"e8"),
  3508 => (x"b1",x"72",x"32",x"c8"),
  3509 => (x"66",x"97",x"e9",x"c0"),
  3510 => (x"b5",x"71",x"4d",x"4a"),
  3511 => (x"c0",x"87",x"f9",x"c0"),
  3512 => (x"49",x"66",x"97",x"e8"),
  3513 => (x"70",x"87",x"f4",x"e5"),
  3514 => (x"eb",x"c0",x"1e",x"49"),
  3515 => (x"e5",x"49",x"66",x"97"),
  3516 => (x"49",x"70",x"87",x"e9"),
  3517 => (x"97",x"ee",x"c0",x"1e"),
  3518 => (x"de",x"e5",x"49",x"66"),
  3519 => (x"49",x"4a",x"70",x"87"),
  3520 => (x"87",x"cb",x"c5",x"ff"),
  3521 => (x"4d",x"70",x"86",x"c8"),
  3522 => (x"c0",x"87",x"cd",x"c0"),
  3523 => (x"49",x"66",x"97",x"e6"),
  3524 => (x"c4",x"87",x"e0",x"e5"),
  3525 => (x"4d",x"bf",x"da",x"cb"),
  3526 => (x"48",x"ca",x"f1",x"c4"),
  3527 => (x"f1",x"c4",x"78",x"c0"),
  3528 => (x"49",x"75",x"5d",x"e3"),
  3529 => (x"c4",x"87",x"c3",x"e2"),
  3530 => (x"c4",x"58",x"df",x"f1"),
  3531 => (x"c4",x"5d",x"f7",x"f1"),
  3532 => (x"c4",x"48",x"f7",x"f1"),
  3533 => (x"78",x"bf",x"ca",x"cb"),
  3534 => (x"48",x"ff",x"f1",x"c4"),
  3535 => (x"66",x"97",x"e5",x"c0"),
  3536 => (x"fb",x"f1",x"c4",x"50"),
  3537 => (x"c4",x"78",x"c1",x"48"),
  3538 => (x"bf",x"97",x"ff",x"f1"),
  3539 => (x"c0",x"05",x"99",x"49"),
  3540 => (x"f1",x"c4",x"87",x"c9"),
  3541 => (x"50",x"c4",x"48",x"ce"),
  3542 => (x"c4",x"87",x"c6",x"c0"),
  3543 => (x"c3",x"48",x"ce",x"f1"),
  3544 => (x"e5",x"49",x"c0",x"50"),
  3545 => (x"e8",x"c8",x"87",x"ed"),
  3546 => (x"87",x"cd",x"e9",x"87"),
  3547 => (x"c8",x"02",x"98",x"70"),
  3548 => (x"ed",x"c0",x"87",x"df"),
  3549 => (x"48",x"49",x"66",x"97"),
  3550 => (x"c0",x"98",x"c0",x"c3"),
  3551 => (x"70",x"58",x"a6",x"e4"),
  3552 => (x"dc",x"c0",x"02",x"98"),
  3553 => (x"c0",x"c1",x"48",x"87"),
  3554 => (x"a6",x"e4",x"c0",x"88"),
  3555 => (x"02",x"98",x"70",x"58"),
  3556 => (x"48",x"87",x"e9",x"c0"),
  3557 => (x"c0",x"88",x"c0",x"c1"),
  3558 => (x"70",x"58",x"a6",x"e4"),
  3559 => (x"c7",x"c1",x"02",x"98"),
  3560 => (x"97",x"e7",x"c0",x"87"),
  3561 => (x"31",x"d0",x"49",x"66"),
  3562 => (x"66",x"97",x"e8",x"c0"),
  3563 => (x"72",x"32",x"c8",x"4a"),
  3564 => (x"97",x"e9",x"c0",x"b1"),
  3565 => (x"71",x"4d",x"4a",x"66"),
  3566 => (x"87",x"ee",x"c1",x"b5"),
  3567 => (x"66",x"97",x"e8",x"c0"),
  3568 => (x"87",x"d7",x"e2",x"49"),
  3569 => (x"c0",x"1e",x"49",x"70"),
  3570 => (x"49",x"66",x"97",x"eb"),
  3571 => (x"70",x"87",x"cc",x"e2"),
  3572 => (x"ee",x"c0",x"1e",x"49"),
  3573 => (x"e2",x"49",x"66",x"97"),
  3574 => (x"4a",x"70",x"87",x"c1"),
  3575 => (x"ee",x"c1",x"ff",x"49"),
  3576 => (x"70",x"86",x"c8",x"87"),
  3577 => (x"87",x"c2",x"c1",x"4d"),
  3578 => (x"66",x"97",x"e6",x"c0"),
  3579 => (x"87",x"eb",x"e1",x"49"),
  3580 => (x"c0",x"48",x"49",x"70"),
  3581 => (x"70",x"58",x"a6",x"e4"),
  3582 => (x"c6",x"c0",x"05",x"98"),
  3583 => (x"a6",x"e0",x"c0",x"87"),
  3584 => (x"c0",x"78",x"c1",x"48"),
  3585 => (x"c4",x"48",x"66",x"e0"),
  3586 => (x"b7",x"bf",x"ce",x"cb"),
  3587 => (x"cc",x"c0",x"06",x"a8"),
  3588 => (x"a6",x"e0",x"c0",x"87"),
  3589 => (x"ca",x"cb",x"c4",x"48"),
  3590 => (x"c9",x"c0",x"78",x"bf"),
  3591 => (x"a6",x"e0",x"c0",x"87"),
  3592 => (x"de",x"cb",x"c4",x"48"),
  3593 => (x"e0",x"c0",x"78",x"bf"),
  3594 => (x"f1",x"c4",x"4d",x"66"),
  3595 => (x"e5",x"c0",x"48",x"ff"),
  3596 => (x"c4",x"50",x"66",x"97"),
  3597 => (x"c4",x"5d",x"fb",x"f1"),
  3598 => (x"bf",x"97",x"ff",x"f1"),
  3599 => (x"c0",x"05",x"99",x"49"),
  3600 => (x"f1",x"c4",x"87",x"c9"),
  3601 => (x"50",x"c0",x"48",x"ce"),
  3602 => (x"c4",x"87",x"c6",x"c0"),
  3603 => (x"c3",x"48",x"ce",x"f1"),
  3604 => (x"ff",x"f1",x"c4",x"50"),
  3605 => (x"c2",x"49",x"bf",x"97"),
  3606 => (x"f4",x"c4",x"02",x"a9"),
  3607 => (x"e1",x"49",x"c0",x"87"),
  3608 => (x"ec",x"c4",x"87",x"cb"),
  3609 => (x"87",x"d1",x"e5",x"87"),
  3610 => (x"c4",x"02",x"98",x"70"),
  3611 => (x"f1",x"c4",x"87",x"e3"),
  3612 => (x"50",x"c4",x"48",x"ce"),
  3613 => (x"f4",x"e0",x"49",x"c0"),
  3614 => (x"87",x"d5",x"c4",x"87"),
  3615 => (x"70",x"87",x"fa",x"e4"),
  3616 => (x"cc",x"c4",x"02",x"98"),
  3617 => (x"df",x"f1",x"c4",x"87"),
  3618 => (x"cb",x"c4",x"48",x"bf"),
  3619 => (x"c0",x"88",x"bf",x"da"),
  3620 => (x"ca",x"58",x"a6",x"e4"),
  3621 => (x"a6",x"c1",x"7e",x"97"),
  3622 => (x"50",x"c0",x"c2",x"48"),
  3623 => (x"97",x"ce",x"f1",x"c4"),
  3624 => (x"f7",x"c0",x"48",x"bf"),
  3625 => (x"a8",x"c4",x"58",x"a6"),
  3626 => (x"87",x"c9",x"c0",x"05"),
  3627 => (x"48",x"a6",x"f3",x"c0"),
  3628 => (x"e1",x"c0",x"78",x"c2"),
  3629 => (x"66",x"f3",x"c0",x"87"),
  3630 => (x"05",x"a8",x"c3",x"48"),
  3631 => (x"c0",x"87",x"c9",x"c0"),
  3632 => (x"c0",x"48",x"a6",x"f7"),
  3633 => (x"87",x"c6",x"c0",x"78"),
  3634 => (x"48",x"a6",x"f7",x"c0"),
  3635 => (x"f3",x"c0",x"78",x"c3"),
  3636 => (x"f7",x"c0",x"48",x"a6"),
  3637 => (x"a6",x"c2",x"78",x"66"),
  3638 => (x"66",x"f3",x"c0",x"48"),
  3639 => (x"c4",x"50",x"c0",x"50"),
  3640 => (x"49",x"bf",x"db",x"f1"),
  3641 => (x"dc",x"ff",x"81",x"c1"),
  3642 => (x"a6",x"c4",x"87",x"fc"),
  3643 => (x"f1",x"c4",x"50",x"08"),
  3644 => (x"ff",x"49",x"bf",x"db"),
  3645 => (x"c5",x"87",x"ef",x"dc"),
  3646 => (x"c0",x"50",x"08",x"a6"),
  3647 => (x"1e",x"4b",x"a6",x"f0"),
  3648 => (x"49",x"66",x"e4",x"c0"),
  3649 => (x"87",x"f7",x"fb",x"fe"),
  3650 => (x"66",x"97",x"f4",x"c0"),
  3651 => (x"d5",x"dc",x"ff",x"49"),
  3652 => (x"08",x"a6",x"ca",x"87"),
  3653 => (x"97",x"f5",x"c0",x"50"),
  3654 => (x"dc",x"ff",x"49",x"66"),
  3655 => (x"a6",x"cb",x"87",x"c8"),
  3656 => (x"f6",x"c0",x"50",x"08"),
  3657 => (x"ff",x"49",x"66",x"97"),
  3658 => (x"cc",x"87",x"fb",x"db"),
  3659 => (x"73",x"50",x"08",x"a6"),
  3660 => (x"df",x"f1",x"c4",x"1e"),
  3661 => (x"fb",x"fe",x"49",x"bf"),
  3662 => (x"f8",x"c0",x"87",x"c5"),
  3663 => (x"ff",x"49",x"66",x"97"),
  3664 => (x"d1",x"87",x"e3",x"db"),
  3665 => (x"c0",x"50",x"08",x"a6"),
  3666 => (x"49",x"66",x"97",x"f9"),
  3667 => (x"87",x"d6",x"db",x"ff"),
  3668 => (x"50",x"08",x"a6",x"d2"),
  3669 => (x"66",x"97",x"fa",x"c0"),
  3670 => (x"c9",x"db",x"ff",x"49"),
  3671 => (x"08",x"a6",x"d3",x"87"),
  3672 => (x"ca",x"1e",x"c1",x"50"),
  3673 => (x"49",x"a6",x"d2",x"1e"),
  3674 => (x"87",x"f5",x"dd",x"ff"),
  3675 => (x"49",x"c0",x"86",x"d0"),
  3676 => (x"87",x"f9",x"dc",x"ff"),
  3677 => (x"c0",x"87",x"da",x"c0"),
  3678 => (x"e0",x"c0",x"1e",x"1e"),
  3679 => (x"ff",x"49",x"c5",x"1e"),
  3680 => (x"cc",x"87",x"d5",x"dc"),
  3681 => (x"d4",x"f1",x"c4",x"86"),
  3682 => (x"c1",x"78",x"c0",x"48"),
  3683 => (x"dc",x"dc",x"ff",x"49"),
  3684 => (x"8e",x"c4",x"ff",x"87"),
  3685 => (x"87",x"fb",x"da",x"ff"),
  3686 => (x"ff",x"86",x"f4",x"1e"),
  3687 => (x"c5",x"c8",x"48",x"d0"),
  3688 => (x"48",x"d4",x"ff",x"78"),
  3689 => (x"c0",x"78",x"e3",x"c1"),
  3690 => (x"48",x"d4",x"ff",x"4a"),
  3691 => (x"49",x"76",x"78",x"c0"),
  3692 => (x"51",x"68",x"81",x"72"),
  3693 => (x"b7",x"ca",x"82",x"c1"),
  3694 => (x"87",x"ed",x"04",x"aa"),
  3695 => (x"c4",x"48",x"d0",x"ff"),
  3696 => (x"26",x"8e",x"f4",x"78"),
  3697 => (x"f1",x"c4",x"1e",x"4f"),
  3698 => (x"50",x"c1",x"48",x"d9"),
  3699 => (x"c4",x"1e",x"4f",x"26"),
  3700 => (x"c0",x"48",x"ca",x"f1"),
  3701 => (x"db",x"f1",x"c4",x"78"),
  3702 => (x"78",x"40",x"c0",x"48"),
  3703 => (x"48",x"e7",x"f1",x"c4"),
  3704 => (x"f1",x"c4",x"78",x"c0"),
  3705 => (x"50",x"c1",x"48",x"cf"),
  3706 => (x"bf",x"f6",x"cb",x"c4"),
  3707 => (x"c0",x"87",x"c4",x"02"),
  3708 => (x"c1",x"87",x"c2",x"49"),
  3709 => (x"d2",x"f1",x"c4",x"49"),
  3710 => (x"f1",x"c4",x"59",x"97"),
  3711 => (x"40",x"c0",x"48",x"eb"),
  3712 => (x"d4",x"f1",x"c4",x"78"),
  3713 => (x"50",x"40",x"c0",x"48"),
  3714 => (x"f3",x"f1",x"c4",x"50"),
  3715 => (x"78",x"40",x"c0",x"48"),
  3716 => (x"48",x"ff",x"f1",x"c4"),
  3717 => (x"78",x"9f",x"50",x"c0"),
  3718 => (x"48",x"da",x"f1",x"c4"),
  3719 => (x"4f",x"26",x"50",x"c1"),
  3720 => (x"ff",x"1e",x"73",x"1e"),
  3721 => (x"c5",x"c8",x"48",x"d0"),
  3722 => (x"48",x"d4",x"ff",x"78"),
  3723 => (x"68",x"78",x"e0",x"c1"),
  3724 => (x"99",x"ff",x"c3",x"49"),
  3725 => (x"c4",x"48",x"d0",x"ff"),
  3726 => (x"49",x"4b",x"71",x"78"),
  3727 => (x"c3",x"02",x"99",x"c1"),
  3728 => (x"87",x"df",x"e6",x"87"),
  3729 => (x"99",x"c2",x"49",x"73"),
  3730 => (x"fd",x"87",x"c3",x"02"),
  3731 => (x"49",x"73",x"87",x"ca"),
  3732 => (x"c3",x"02",x"99",x"c4"),
  3733 => (x"87",x"ed",x"fd",x"87"),
  3734 => (x"99",x"c8",x"49",x"73"),
  3735 => (x"fd",x"87",x"d6",x"02"),
  3736 => (x"d0",x"ff",x"87",x"ec"),
  3737 => (x"78",x"c5",x"c8",x"48"),
  3738 => (x"c1",x"48",x"d4",x"ff"),
  3739 => (x"78",x"c0",x"78",x"e6"),
  3740 => (x"c4",x"48",x"d0",x"ff"),
  3741 => (x"d0",x"49",x"73",x"78"),
  3742 => (x"de",x"f1",x"c4",x"99"),
  3743 => (x"dd",x"ff",x"59",x"97"),
  3744 => (x"f1",x"c4",x"87",x"de"),
  3745 => (x"d7",x"02",x"bf",x"d4"),
  3746 => (x"ca",x"f1",x"c4",x"87"),
  3747 => (x"87",x"d0",x"05",x"bf"),
  3748 => (x"9f",x"c0",x"f2",x"c4"),
  3749 => (x"d8",x"ff",x"49",x"bf"),
  3750 => (x"f1",x"c4",x"87",x"d3"),
  3751 => (x"78",x"c0",x"48",x"d4"),
  3752 => (x"97",x"d8",x"f1",x"c4"),
  3753 => (x"87",x"d9",x"02",x"bf"),
  3754 => (x"c8",x"48",x"d0",x"ff"),
  3755 => (x"d4",x"ff",x"78",x"c5"),
  3756 => (x"78",x"e5",x"c1",x"48"),
  3757 => (x"d0",x"ff",x"78",x"c0"),
  3758 => (x"c4",x"78",x"c4",x"48"),
  3759 => (x"c0",x"48",x"d8",x"f1"),
  3760 => (x"d2",x"d6",x"ff",x"50"),
  3761 => (x"00",x"00",x"00",x"87"),
  3762 => (x"4a",x"71",x"1e",x"00"),
  3763 => (x"49",x"bf",x"c8",x"ff"),
  3764 => (x"26",x"48",x"a1",x"72"),
  3765 => (x"c8",x"ff",x"1e",x"4f"),
  3766 => (x"c0",x"fe",x"89",x"bf"),
  3767 => (x"c0",x"c0",x"c0",x"c0"),
  3768 => (x"87",x"c4",x"01",x"a9"),
  3769 => (x"87",x"c2",x"4a",x"c0"),
  3770 => (x"48",x"72",x"4a",x"c1"),
  3771 => (x"5e",x"0e",x"4f",x"26"),
  3772 => (x"0e",x"5d",x"5c",x"5b"),
  3773 => (x"d4",x"ff",x"4b",x"71"),
  3774 => (x"48",x"66",x"d0",x"4c"),
  3775 => (x"49",x"d6",x"78",x"c0"),
  3776 => (x"87",x"df",x"cf",x"fe"),
  3777 => (x"6c",x"7c",x"ff",x"c3"),
  3778 => (x"99",x"ff",x"c3",x"49"),
  3779 => (x"c3",x"49",x"4d",x"71"),
  3780 => (x"e0",x"c1",x"99",x"f0"),
  3781 => (x"87",x"cb",x"05",x"a9"),
  3782 => (x"6c",x"7c",x"ff",x"c3"),
  3783 => (x"d0",x"98",x"c3",x"48"),
  3784 => (x"c3",x"78",x"08",x"66"),
  3785 => (x"4a",x"6c",x"7c",x"ff"),
  3786 => (x"c3",x"31",x"c8",x"49"),
  3787 => (x"4a",x"6c",x"7c",x"ff"),
  3788 => (x"49",x"72",x"b2",x"71"),
  3789 => (x"ff",x"c3",x"31",x"c8"),
  3790 => (x"71",x"4a",x"6c",x"7c"),
  3791 => (x"c8",x"49",x"72",x"b2"),
  3792 => (x"7c",x"ff",x"c3",x"31"),
  3793 => (x"b2",x"71",x"4a",x"6c"),
  3794 => (x"c0",x"48",x"d0",x"ff"),
  3795 => (x"9b",x"73",x"78",x"e0"),
  3796 => (x"72",x"87",x"c2",x"02"),
  3797 => (x"26",x"48",x"75",x"7b"),
  3798 => (x"26",x"4c",x"26",x"4d"),
  3799 => (x"1e",x"4f",x"26",x"4b"),
  3800 => (x"5e",x"0e",x"4f",x"26"),
  3801 => (x"f8",x"0e",x"5c",x"5b"),
  3802 => (x"c8",x"1e",x"76",x"86"),
  3803 => (x"fd",x"fd",x"49",x"a6"),
  3804 => (x"70",x"86",x"c4",x"87"),
  3805 => (x"c0",x"48",x"6e",x"4b"),
  3806 => (x"f0",x"c2",x"01",x"a8"),
  3807 => (x"c3",x"4a",x"73",x"87"),
  3808 => (x"d0",x"c1",x"9a",x"f0"),
  3809 => (x"87",x"c7",x"02",x"aa"),
  3810 => (x"05",x"aa",x"e0",x"c1"),
  3811 => (x"73",x"87",x"de",x"c2"),
  3812 => (x"02",x"99",x"c8",x"49"),
  3813 => (x"c6",x"ff",x"87",x"c3"),
  3814 => (x"c3",x"4c",x"73",x"87"),
  3815 => (x"05",x"ac",x"c2",x"9c"),
  3816 => (x"c4",x"87",x"c2",x"c1"),
  3817 => (x"31",x"c9",x"49",x"66"),
  3818 => (x"66",x"c4",x"1e",x"71"),
  3819 => (x"c4",x"92",x"d4",x"4a"),
  3820 => (x"72",x"49",x"c2",x"f2"),
  3821 => (x"f7",x"fe",x"fc",x"81"),
  3822 => (x"fe",x"49",x"d8",x"87"),
  3823 => (x"c8",x"87",x"e4",x"cc"),
  3824 => (x"f9",x"c3",x"1e",x"c0"),
  3825 => (x"db",x"fc",x"49",x"fa"),
  3826 => (x"d0",x"ff",x"87",x"d0"),
  3827 => (x"78",x"e0",x"c0",x"48"),
  3828 => (x"1e",x"fa",x"f9",x"c3"),
  3829 => (x"d4",x"4a",x"66",x"cc"),
  3830 => (x"c2",x"f2",x"c4",x"92"),
  3831 => (x"fc",x"81",x"72",x"49"),
  3832 => (x"cc",x"87",x"ca",x"fd"),
  3833 => (x"05",x"ac",x"c1",x"86"),
  3834 => (x"c4",x"87",x"c2",x"c1"),
  3835 => (x"31",x"c9",x"49",x"66"),
  3836 => (x"66",x"c4",x"1e",x"71"),
  3837 => (x"c4",x"92",x"d4",x"4a"),
  3838 => (x"72",x"49",x"c2",x"f2"),
  3839 => (x"ef",x"fd",x"fc",x"81"),
  3840 => (x"fa",x"f9",x"c3",x"87"),
  3841 => (x"4a",x"66",x"c8",x"1e"),
  3842 => (x"f2",x"c4",x"92",x"d4"),
  3843 => (x"81",x"72",x"49",x"c2"),
  3844 => (x"87",x"d6",x"fb",x"fc"),
  3845 => (x"cb",x"fe",x"49",x"d7"),
  3846 => (x"c0",x"c8",x"87",x"c9"),
  3847 => (x"fa",x"f9",x"c3",x"1e"),
  3848 => (x"df",x"d9",x"fc",x"49"),
  3849 => (x"ff",x"86",x"cc",x"87"),
  3850 => (x"e0",x"c0",x"48",x"d0"),
  3851 => (x"fc",x"8e",x"f8",x"78"),
  3852 => (x"5e",x"0e",x"87",x"e7"),
  3853 => (x"0e",x"5d",x"5c",x"5b"),
  3854 => (x"ff",x"4d",x"71",x"1e"),
  3855 => (x"66",x"d4",x"4c",x"d4"),
  3856 => (x"b7",x"c3",x"48",x"7e"),
  3857 => (x"87",x"c5",x"06",x"a8"),
  3858 => (x"e2",x"c1",x"48",x"c0"),
  3859 => (x"fd",x"49",x"75",x"87"),
  3860 => (x"75",x"87",x"db",x"d1"),
  3861 => (x"4b",x"66",x"c4",x"1e"),
  3862 => (x"f2",x"c4",x"93",x"d4"),
  3863 => (x"49",x"73",x"83",x"c2"),
  3864 => (x"87",x"ea",x"f6",x"fc"),
  3865 => (x"4b",x"6b",x"83",x"c8"),
  3866 => (x"c8",x"48",x"d0",x"ff"),
  3867 => (x"7c",x"dd",x"78",x"e1"),
  3868 => (x"ff",x"c3",x"49",x"73"),
  3869 => (x"73",x"7c",x"71",x"99"),
  3870 => (x"29",x"b7",x"c8",x"49"),
  3871 => (x"71",x"99",x"ff",x"c3"),
  3872 => (x"d0",x"49",x"73",x"7c"),
  3873 => (x"ff",x"c3",x"29",x"b7"),
  3874 => (x"73",x"7c",x"71",x"99"),
  3875 => (x"29",x"b7",x"d8",x"49"),
  3876 => (x"7c",x"c0",x"7c",x"71"),
  3877 => (x"7c",x"7c",x"7c",x"7c"),
  3878 => (x"7c",x"7c",x"7c",x"7c"),
  3879 => (x"c0",x"7c",x"7c",x"7c"),
  3880 => (x"66",x"c4",x"78",x"e0"),
  3881 => (x"fe",x"49",x"dc",x"1e"),
  3882 => (x"c8",x"87",x"dd",x"c9"),
  3883 => (x"26",x"48",x"73",x"86"),
  3884 => (x"0e",x"87",x"e4",x"fa"),
  3885 => (x"5d",x"5c",x"5b",x"5e"),
  3886 => (x"7e",x"71",x"1e",x"0e"),
  3887 => (x"6e",x"4b",x"d4",x"ff"),
  3888 => (x"d6",x"f2",x"c4",x"1e"),
  3889 => (x"c5",x"f5",x"fc",x"49"),
  3890 => (x"70",x"86",x"c4",x"87"),
  3891 => (x"c3",x"02",x"9d",x"4d"),
  3892 => (x"f2",x"c4",x"87",x"c3"),
  3893 => (x"6e",x"4c",x"bf",x"de"),
  3894 => (x"d1",x"cf",x"fd",x"49"),
  3895 => (x"48",x"d0",x"ff",x"87"),
  3896 => (x"c1",x"78",x"c5",x"c8"),
  3897 => (x"4a",x"c0",x"7b",x"d6"),
  3898 => (x"82",x"c1",x"7b",x"15"),
  3899 => (x"aa",x"b7",x"e0",x"c0"),
  3900 => (x"ff",x"87",x"f5",x"04"),
  3901 => (x"78",x"c4",x"48",x"d0"),
  3902 => (x"c1",x"78",x"c5",x"c8"),
  3903 => (x"7b",x"c1",x"7b",x"d3"),
  3904 => (x"9c",x"74",x"78",x"c4"),
  3905 => (x"87",x"fc",x"c1",x"02"),
  3906 => (x"7e",x"fa",x"f9",x"c3"),
  3907 => (x"8c",x"4d",x"c0",x"c8"),
  3908 => (x"03",x"ac",x"b7",x"c0"),
  3909 => (x"c0",x"c8",x"87",x"c6"),
  3910 => (x"4c",x"c0",x"4d",x"a4"),
  3911 => (x"97",x"eb",x"c6",x"c4"),
  3912 => (x"99",x"d0",x"49",x"bf"),
  3913 => (x"c0",x"87",x"d2",x"02"),
  3914 => (x"d6",x"f2",x"c4",x"1e"),
  3915 => (x"f9",x"f6",x"fc",x"49"),
  3916 => (x"70",x"86",x"c4",x"87"),
  3917 => (x"ef",x"c0",x"4a",x"49"),
  3918 => (x"fa",x"f9",x"c3",x"87"),
  3919 => (x"d6",x"f2",x"c4",x"1e"),
  3920 => (x"e5",x"f6",x"fc",x"49"),
  3921 => (x"70",x"86",x"c4",x"87"),
  3922 => (x"d0",x"ff",x"4a",x"49"),
  3923 => (x"78",x"c5",x"c8",x"48"),
  3924 => (x"6e",x"7b",x"d4",x"c1"),
  3925 => (x"6e",x"7b",x"bf",x"97"),
  3926 => (x"70",x"80",x"c1",x"48"),
  3927 => (x"05",x"8d",x"c1",x"7e"),
  3928 => (x"ff",x"87",x"f0",x"ff"),
  3929 => (x"78",x"c4",x"48",x"d0"),
  3930 => (x"c5",x"05",x"9a",x"72"),
  3931 => (x"c0",x"48",x"c0",x"87"),
  3932 => (x"1e",x"c1",x"87",x"e5"),
  3933 => (x"49",x"d6",x"f2",x"c4"),
  3934 => (x"87",x"cd",x"f4",x"fc"),
  3935 => (x"9c",x"74",x"86",x"c4"),
  3936 => (x"87",x"c4",x"fe",x"05"),
  3937 => (x"c8",x"48",x"d0",x"ff"),
  3938 => (x"d3",x"c1",x"78",x"c5"),
  3939 => (x"c4",x"7b",x"c0",x"7b"),
  3940 => (x"c2",x"48",x"c1",x"78"),
  3941 => (x"26",x"48",x"c0",x"87"),
  3942 => (x"4c",x"26",x"4d",x"26"),
  3943 => (x"4f",x"26",x"4b",x"26"),
  3944 => (x"5c",x"5b",x"5e",x"0e"),
  3945 => (x"cc",x"4b",x"71",x"0e"),
  3946 => (x"87",x"dd",x"02",x"66"),
  3947 => (x"8c",x"f0",x"c0",x"4c"),
  3948 => (x"74",x"87",x"dd",x"02"),
  3949 => (x"02",x"8a",x"c1",x"4a"),
  3950 => (x"02",x"8a",x"87",x"d6"),
  3951 => (x"02",x"8a",x"87",x"d2"),
  3952 => (x"8a",x"d0",x"87",x"ce"),
  3953 => (x"df",x"87",x"db",x"02"),
  3954 => (x"fb",x"49",x"73",x"87"),
  3955 => (x"87",x"d8",x"87",x"e5"),
  3956 => (x"49",x"c0",x"1e",x"74"),
  3957 => (x"74",x"87",x"db",x"f9"),
  3958 => (x"f9",x"49",x"73",x"1e"),
  3959 => (x"86",x"c8",x"87",x"d4"),
  3960 => (x"49",x"73",x"87",x"c6"),
  3961 => (x"87",x"dd",x"d0",x"fd"),
  3962 => (x"00",x"87",x"ef",x"fe"),
  3963 => (x"fa",x"f8",x"c3",x"1e"),
  3964 => (x"b9",x"c1",x"49",x"bf"),
  3965 => (x"59",x"fe",x"f8",x"c3"),
  3966 => (x"c3",x"48",x"d4",x"ff"),
  3967 => (x"d0",x"ff",x"78",x"ff"),
  3968 => (x"78",x"e1",x"c8",x"48"),
  3969 => (x"c1",x"48",x"d4",x"ff"),
  3970 => (x"71",x"31",x"c4",x"78"),
  3971 => (x"48",x"d0",x"ff",x"78"),
  3972 => (x"26",x"78",x"e0",x"c0"),
  3973 => (x"f8",x"c3",x"1e",x"4f"),
  3974 => (x"f2",x"c4",x"1e",x"ee"),
  3975 => (x"ef",x"fc",x"49",x"d6"),
  3976 => (x"86",x"c4",x"87",x"ec"),
  3977 => (x"c3",x"02",x"98",x"70"),
  3978 => (x"87",x"c0",x"ff",x"87"),
  3979 => (x"35",x"31",x"4f",x"26"),
  3980 => (x"20",x"5a",x"48",x"4b"),
  3981 => (x"46",x"43",x"20",x"20"),
  3982 => (x"00",x"00",x"00",x"47"),
  3983 => (x"9f",x"1a",x"00",x"00"),
  3984 => (x"14",x"11",x"12",x"58"),
  3985 => (x"23",x"1c",x"1b",x"1d"),
  3986 => (x"59",x"5a",x"a7",x"4a"),
  3987 => (x"f2",x"f5",x"94",x"91"),
  3988 => (x"f2",x"f5",x"f4",x"eb"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

